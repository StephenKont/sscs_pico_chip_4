magic
tech sky130A
magscale 1 2
timestamp 1666550119
<< metal3 >>
rect -2663 7300 -2381 7456
rect 2251 7300 2543 7448
rect -4909 5304 -147 7300
rect 17 5304 4909 7300
rect -4909 4876 4909 5304
rect -4909 2612 -147 4876
rect -4909 2500 -173 2612
rect 17 2500 4909 4876
rect -2663 2400 -2381 2500
rect 2251 2400 2543 2500
rect -4909 24 -173 2400
rect 15 24 4909 2400
rect -4909 -404 4909 24
rect -4909 -2400 -173 -404
rect 15 -2400 4909 -404
rect -2663 -2500 -2381 -2400
rect 2251 -2500 2543 -2400
rect -4909 -4812 -173 -2500
rect 15 -4812 4909 -2500
rect -4909 -5240 4909 -4812
rect -4909 -7300 -173 -5240
rect 15 -7300 4909 -5240
rect -2663 -7390 -2381 -7300
rect 2251 -7450 2543 -7300
<< mimcap >>
rect -4809 7160 -209 7200
rect -4809 2640 -4769 7160
rect -249 2640 -209 7160
rect -4809 2600 -209 2640
rect 110 7160 4710 7200
rect 110 2640 150 7160
rect 4670 2640 4710 7160
rect 110 2600 4710 2640
rect -4809 2260 -209 2300
rect -4809 -2260 -4769 2260
rect -249 -2260 -209 2260
rect -4809 -2300 -209 -2260
rect 110 2260 4710 2300
rect 110 -2260 150 2260
rect 4670 -2260 4710 2260
rect 110 -2300 4710 -2260
rect -4809 -2640 -209 -2600
rect -4809 -7160 -4769 -2640
rect -249 -7160 -209 -2640
rect -4809 -7200 -209 -7160
rect 110 -2640 4710 -2600
rect 110 -7160 150 -2640
rect 4670 -7160 4710 -2640
rect 110 -7200 4710 -7160
<< mimcapcontact >>
rect -4769 2640 -249 7160
rect 150 2640 4670 7160
rect -4769 -2260 -249 2260
rect 150 -2260 4670 2260
rect -4769 -7160 -249 -2640
rect 150 -7160 4670 -2640
<< metal4 >>
rect -2607 7161 -2411 7402
rect 2297 7161 2507 7408
rect -4770 7160 -248 7161
rect -4770 2640 -4769 7160
rect -249 5298 -248 7160
rect 149 7160 4671 7161
rect 149 5298 150 7160
rect -249 4870 150 5298
rect -249 2640 -248 4870
rect -4770 2639 -248 2640
rect 149 2640 150 4870
rect 4670 2640 4671 7160
rect 149 2639 4671 2640
rect -2607 2261 -2411 2639
rect 2297 2261 2507 2639
rect -4770 2260 -248 2261
rect -4770 -2260 -4769 2260
rect -249 14 -248 2260
rect 149 2260 4671 2261
rect 149 14 150 2260
rect -249 -414 150 14
rect -249 -2260 -248 -414
rect -4770 -2261 -248 -2260
rect 149 -2260 150 -414
rect 4670 -2260 4671 2260
rect 149 -2261 4671 -2260
rect -2607 -2639 -2411 -2261
rect 2297 -2639 2507 -2261
rect -4770 -2640 -248 -2639
rect -4770 -7160 -4769 -2640
rect -249 -4808 -248 -2640
rect 149 -2640 4671 -2639
rect 149 -4808 150 -2640
rect -249 -5236 150 -4808
rect -249 -7160 -248 -5236
rect -4770 -7161 -248 -7160
rect 149 -7160 150 -5236
rect 4670 -7160 4671 -2640
rect 149 -7161 4671 -7160
rect -2607 -7332 -2411 -7161
rect -2561 -7350 -2457 -7332
rect 2297 -7426 2507 -7161
use sky130_fd_pr__cap_mim_m3_2_3VRXMH  sky130_fd_pr__cap_mim_m3_2_3VRXMH_0
timestamp 1666550119
transform 1 0 521 0 1 32
box -5312 -7364 5004 7384
<< properties >>
string FIXED_BBOX 10 2500 4810 7300
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 23.00 l 23.00 val 1.075k carea 2.00 cperi 0.19 nx 2 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
