magic
tech sky130A
magscale 1 2
timestamp 1668293870
<< pwell >>
rect -475 -1210 475 1210
<< nmos >>
rect -279 -1000 -29 1000
rect 29 -1000 279 1000
<< ndiff >>
rect -337 988 -279 1000
rect -337 -988 -325 988
rect -291 -988 -279 988
rect -337 -1000 -279 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 279 988 337 1000
rect 279 -988 291 988
rect 325 -988 337 988
rect 279 -1000 337 -988
<< ndiffc >>
rect -325 -988 -291 988
rect -17 -988 17 988
rect 291 -988 325 988
<< psubdiff >>
rect -439 1140 -343 1174
rect 343 1140 439 1174
rect -439 1078 -405 1140
rect 405 1078 439 1140
rect -439 -1140 -405 -1078
rect 405 -1140 439 -1078
rect -439 -1174 -343 -1140
rect 343 -1174 439 -1140
<< psubdiffcont >>
rect -343 1140 343 1174
rect -439 -1078 -405 1078
rect 405 -1078 439 1078
rect -343 -1174 343 -1140
<< poly >>
rect -279 1072 -29 1088
rect -279 1038 -263 1072
rect -45 1038 -29 1072
rect -279 1000 -29 1038
rect 29 1072 279 1088
rect 29 1038 45 1072
rect 263 1038 279 1072
rect 29 1000 279 1038
rect -279 -1038 -29 -1000
rect -279 -1072 -263 -1038
rect -45 -1072 -29 -1038
rect -279 -1088 -29 -1072
rect 29 -1038 279 -1000
rect 29 -1072 45 -1038
rect 263 -1072 279 -1038
rect 29 -1088 279 -1072
<< polycont >>
rect -263 1038 -45 1072
rect 45 1038 263 1072
rect -263 -1072 -45 -1038
rect 45 -1072 263 -1038
<< locali >>
rect -439 1140 -343 1174
rect 343 1140 439 1174
rect -439 1078 -405 1140
rect 405 1078 439 1140
rect -279 1038 -263 1072
rect -45 1038 -29 1072
rect 29 1038 45 1072
rect 263 1038 279 1072
rect -325 988 -291 1004
rect -325 -1004 -291 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 291 988 325 1004
rect 291 -1004 325 -988
rect -279 -1072 -263 -1038
rect -45 -1072 -29 -1038
rect 29 -1072 45 -1038
rect 263 -1072 279 -1038
rect -439 -1140 -405 -1078
rect 405 -1140 439 -1078
rect -439 -1174 -343 -1140
rect 343 -1174 439 -1140
<< viali >>
rect -263 1038 -45 1072
rect 45 1038 263 1072
rect -325 -988 -291 988
rect -17 -988 17 988
rect 291 -988 325 988
rect -263 -1072 -45 -1038
rect 45 -1072 263 -1038
<< metal1 >>
rect -275 1072 -33 1078
rect -275 1038 -263 1072
rect -45 1038 -33 1072
rect -275 1032 -33 1038
rect 33 1072 275 1078
rect 33 1038 45 1072
rect 263 1038 275 1072
rect 33 1032 275 1038
rect -331 988 -285 1000
rect -331 -988 -325 988
rect -291 -988 -285 988
rect -331 -1000 -285 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 285 988 331 1000
rect 285 -988 291 988
rect 325 -988 331 988
rect 285 -1000 331 -988
rect -275 -1038 -33 -1032
rect -275 -1072 -263 -1038
rect -45 -1072 -33 -1038
rect -275 -1078 -33 -1072
rect 33 -1038 275 -1032
rect 33 -1072 45 -1038
rect 263 -1072 275 -1038
rect 33 -1078 275 -1072
<< properties >>
string FIXED_BBOX -422 -1157 422 1157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 1.25 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
