magic
tech sky130A
magscale 1 2
timestamp 1665420977
<< nwell >>
rect -308 -2857 308 2857
<< mvpmos >>
rect -50 2360 50 2560
rect -50 2032 50 2232
rect -50 1704 50 1904
rect -50 1376 50 1576
rect -50 1048 50 1248
rect -50 720 50 920
rect -50 392 50 592
rect -50 64 50 264
rect -50 -264 50 -64
rect -50 -592 50 -392
rect -50 -920 50 -720
rect -50 -1248 50 -1048
rect -50 -1576 50 -1376
rect -50 -1904 50 -1704
rect -50 -2232 50 -2032
rect -50 -2560 50 -2360
<< mvpdiff >>
rect -108 2548 -50 2560
rect -108 2372 -96 2548
rect -62 2372 -50 2548
rect -108 2360 -50 2372
rect 50 2548 108 2560
rect 50 2372 62 2548
rect 96 2372 108 2548
rect 50 2360 108 2372
rect -108 2220 -50 2232
rect -108 2044 -96 2220
rect -62 2044 -50 2220
rect -108 2032 -50 2044
rect 50 2220 108 2232
rect 50 2044 62 2220
rect 96 2044 108 2220
rect 50 2032 108 2044
rect -108 1892 -50 1904
rect -108 1716 -96 1892
rect -62 1716 -50 1892
rect -108 1704 -50 1716
rect 50 1892 108 1904
rect 50 1716 62 1892
rect 96 1716 108 1892
rect 50 1704 108 1716
rect -108 1564 -50 1576
rect -108 1388 -96 1564
rect -62 1388 -50 1564
rect -108 1376 -50 1388
rect 50 1564 108 1576
rect 50 1388 62 1564
rect 96 1388 108 1564
rect 50 1376 108 1388
rect -108 1236 -50 1248
rect -108 1060 -96 1236
rect -62 1060 -50 1236
rect -108 1048 -50 1060
rect 50 1236 108 1248
rect 50 1060 62 1236
rect 96 1060 108 1236
rect 50 1048 108 1060
rect -108 908 -50 920
rect -108 732 -96 908
rect -62 732 -50 908
rect -108 720 -50 732
rect 50 908 108 920
rect 50 732 62 908
rect 96 732 108 908
rect 50 720 108 732
rect -108 580 -50 592
rect -108 404 -96 580
rect -62 404 -50 580
rect -108 392 -50 404
rect 50 580 108 592
rect 50 404 62 580
rect 96 404 108 580
rect 50 392 108 404
rect -108 252 -50 264
rect -108 76 -96 252
rect -62 76 -50 252
rect -108 64 -50 76
rect 50 252 108 264
rect 50 76 62 252
rect 96 76 108 252
rect 50 64 108 76
rect -108 -76 -50 -64
rect -108 -252 -96 -76
rect -62 -252 -50 -76
rect -108 -264 -50 -252
rect 50 -76 108 -64
rect 50 -252 62 -76
rect 96 -252 108 -76
rect 50 -264 108 -252
rect -108 -404 -50 -392
rect -108 -580 -96 -404
rect -62 -580 -50 -404
rect -108 -592 -50 -580
rect 50 -404 108 -392
rect 50 -580 62 -404
rect 96 -580 108 -404
rect 50 -592 108 -580
rect -108 -732 -50 -720
rect -108 -908 -96 -732
rect -62 -908 -50 -732
rect -108 -920 -50 -908
rect 50 -732 108 -720
rect 50 -908 62 -732
rect 96 -908 108 -732
rect 50 -920 108 -908
rect -108 -1060 -50 -1048
rect -108 -1236 -96 -1060
rect -62 -1236 -50 -1060
rect -108 -1248 -50 -1236
rect 50 -1060 108 -1048
rect 50 -1236 62 -1060
rect 96 -1236 108 -1060
rect 50 -1248 108 -1236
rect -108 -1388 -50 -1376
rect -108 -1564 -96 -1388
rect -62 -1564 -50 -1388
rect -108 -1576 -50 -1564
rect 50 -1388 108 -1376
rect 50 -1564 62 -1388
rect 96 -1564 108 -1388
rect 50 -1576 108 -1564
rect -108 -1716 -50 -1704
rect -108 -1892 -96 -1716
rect -62 -1892 -50 -1716
rect -108 -1904 -50 -1892
rect 50 -1716 108 -1704
rect 50 -1892 62 -1716
rect 96 -1892 108 -1716
rect 50 -1904 108 -1892
rect -108 -2044 -50 -2032
rect -108 -2220 -96 -2044
rect -62 -2220 -50 -2044
rect -108 -2232 -50 -2220
rect 50 -2044 108 -2032
rect 50 -2220 62 -2044
rect 96 -2220 108 -2044
rect 50 -2232 108 -2220
rect -108 -2372 -50 -2360
rect -108 -2548 -96 -2372
rect -62 -2548 -50 -2372
rect -108 -2560 -50 -2548
rect 50 -2372 108 -2360
rect 50 -2548 62 -2372
rect 96 -2548 108 -2372
rect 50 -2560 108 -2548
<< mvpdiffc >>
rect -96 2372 -62 2548
rect 62 2372 96 2548
rect -96 2044 -62 2220
rect 62 2044 96 2220
rect -96 1716 -62 1892
rect 62 1716 96 1892
rect -96 1388 -62 1564
rect 62 1388 96 1564
rect -96 1060 -62 1236
rect 62 1060 96 1236
rect -96 732 -62 908
rect 62 732 96 908
rect -96 404 -62 580
rect 62 404 96 580
rect -96 76 -62 252
rect 62 76 96 252
rect -96 -252 -62 -76
rect 62 -252 96 -76
rect -96 -580 -62 -404
rect 62 -580 96 -404
rect -96 -908 -62 -732
rect 62 -908 96 -732
rect -96 -1236 -62 -1060
rect 62 -1236 96 -1060
rect -96 -1564 -62 -1388
rect 62 -1564 96 -1388
rect -96 -1892 -62 -1716
rect 62 -1892 96 -1716
rect -96 -2220 -62 -2044
rect 62 -2220 96 -2044
rect -96 -2548 -62 -2372
rect 62 -2548 96 -2372
<< mvnsubdiff >>
rect -242 2779 242 2791
rect -242 2745 -134 2779
rect 134 2745 242 2779
rect -242 2733 242 2745
rect -242 2683 -184 2733
rect -242 -2683 -230 2683
rect -196 -2683 -184 2683
rect 184 2683 242 2733
rect -242 -2733 -184 -2683
rect 184 -2683 196 2683
rect 230 -2683 242 2683
rect 184 -2733 242 -2683
rect -242 -2745 242 -2733
rect -242 -2779 -134 -2745
rect 134 -2779 242 -2745
rect -242 -2791 242 -2779
<< mvnsubdiffcont >>
rect -134 2745 134 2779
rect -230 -2683 -196 2683
rect 196 -2683 230 2683
rect -134 -2779 134 -2745
<< poly >>
rect -50 2641 50 2657
rect -50 2607 -34 2641
rect 34 2607 50 2641
rect -50 2560 50 2607
rect -50 2313 50 2360
rect -50 2279 -34 2313
rect 34 2279 50 2313
rect -50 2232 50 2279
rect -50 1985 50 2032
rect -50 1951 -34 1985
rect 34 1951 50 1985
rect -50 1904 50 1951
rect -50 1657 50 1704
rect -50 1623 -34 1657
rect 34 1623 50 1657
rect -50 1576 50 1623
rect -50 1329 50 1376
rect -50 1295 -34 1329
rect 34 1295 50 1329
rect -50 1248 50 1295
rect -50 1001 50 1048
rect -50 967 -34 1001
rect 34 967 50 1001
rect -50 920 50 967
rect -50 673 50 720
rect -50 639 -34 673
rect 34 639 50 673
rect -50 592 50 639
rect -50 345 50 392
rect -50 311 -34 345
rect 34 311 50 345
rect -50 264 50 311
rect -50 17 50 64
rect -50 -17 -34 17
rect 34 -17 50 17
rect -50 -64 50 -17
rect -50 -311 50 -264
rect -50 -345 -34 -311
rect 34 -345 50 -311
rect -50 -392 50 -345
rect -50 -639 50 -592
rect -50 -673 -34 -639
rect 34 -673 50 -639
rect -50 -720 50 -673
rect -50 -967 50 -920
rect -50 -1001 -34 -967
rect 34 -1001 50 -967
rect -50 -1048 50 -1001
rect -50 -1295 50 -1248
rect -50 -1329 -34 -1295
rect 34 -1329 50 -1295
rect -50 -1376 50 -1329
rect -50 -1623 50 -1576
rect -50 -1657 -34 -1623
rect 34 -1657 50 -1623
rect -50 -1704 50 -1657
rect -50 -1951 50 -1904
rect -50 -1985 -34 -1951
rect 34 -1985 50 -1951
rect -50 -2032 50 -1985
rect -50 -2279 50 -2232
rect -50 -2313 -34 -2279
rect 34 -2313 50 -2279
rect -50 -2360 50 -2313
rect -50 -2607 50 -2560
rect -50 -2641 -34 -2607
rect 34 -2641 50 -2607
rect -50 -2657 50 -2641
<< polycont >>
rect -34 2607 34 2641
rect -34 2279 34 2313
rect -34 1951 34 1985
rect -34 1623 34 1657
rect -34 1295 34 1329
rect -34 967 34 1001
rect -34 639 34 673
rect -34 311 34 345
rect -34 -17 34 17
rect -34 -345 34 -311
rect -34 -673 34 -639
rect -34 -1001 34 -967
rect -34 -1329 34 -1295
rect -34 -1657 34 -1623
rect -34 -1985 34 -1951
rect -34 -2313 34 -2279
rect -34 -2641 34 -2607
<< locali >>
rect -230 2745 -134 2779
rect 134 2745 230 2779
rect -230 2683 -196 2745
rect 196 2683 230 2745
rect -50 2607 -34 2641
rect 34 2607 50 2641
rect -96 2548 -62 2564
rect -96 2356 -62 2372
rect 62 2548 96 2564
rect 62 2356 96 2372
rect -50 2279 -34 2313
rect 34 2279 50 2313
rect -96 2220 -62 2236
rect -96 2028 -62 2044
rect 62 2220 96 2236
rect 62 2028 96 2044
rect -50 1951 -34 1985
rect 34 1951 50 1985
rect -96 1892 -62 1908
rect -96 1700 -62 1716
rect 62 1892 96 1908
rect 62 1700 96 1716
rect -50 1623 -34 1657
rect 34 1623 50 1657
rect -96 1564 -62 1580
rect -96 1372 -62 1388
rect 62 1564 96 1580
rect 62 1372 96 1388
rect -50 1295 -34 1329
rect 34 1295 50 1329
rect -96 1236 -62 1252
rect -96 1044 -62 1060
rect 62 1236 96 1252
rect 62 1044 96 1060
rect -50 967 -34 1001
rect 34 967 50 1001
rect -96 908 -62 924
rect -96 716 -62 732
rect 62 908 96 924
rect 62 716 96 732
rect -50 639 -34 673
rect 34 639 50 673
rect -96 580 -62 596
rect -96 388 -62 404
rect 62 580 96 596
rect 62 388 96 404
rect -50 311 -34 345
rect 34 311 50 345
rect -96 252 -62 268
rect -96 60 -62 76
rect 62 252 96 268
rect 62 60 96 76
rect -50 -17 -34 17
rect 34 -17 50 17
rect -96 -76 -62 -60
rect -96 -268 -62 -252
rect 62 -76 96 -60
rect 62 -268 96 -252
rect -50 -345 -34 -311
rect 34 -345 50 -311
rect -96 -404 -62 -388
rect -96 -596 -62 -580
rect 62 -404 96 -388
rect 62 -596 96 -580
rect -50 -673 -34 -639
rect 34 -673 50 -639
rect -96 -732 -62 -716
rect -96 -924 -62 -908
rect 62 -732 96 -716
rect 62 -924 96 -908
rect -50 -1001 -34 -967
rect 34 -1001 50 -967
rect -96 -1060 -62 -1044
rect -96 -1252 -62 -1236
rect 62 -1060 96 -1044
rect 62 -1252 96 -1236
rect -50 -1329 -34 -1295
rect 34 -1329 50 -1295
rect -96 -1388 -62 -1372
rect -96 -1580 -62 -1564
rect 62 -1388 96 -1372
rect 62 -1580 96 -1564
rect -50 -1657 -34 -1623
rect 34 -1657 50 -1623
rect -96 -1716 -62 -1700
rect -96 -1908 -62 -1892
rect 62 -1716 96 -1700
rect 62 -1908 96 -1892
rect -50 -1985 -34 -1951
rect 34 -1985 50 -1951
rect -96 -2044 -62 -2028
rect -96 -2236 -62 -2220
rect 62 -2044 96 -2028
rect 62 -2236 96 -2220
rect -50 -2313 -34 -2279
rect 34 -2313 50 -2279
rect -96 -2372 -62 -2356
rect -96 -2564 -62 -2548
rect 62 -2372 96 -2356
rect 62 -2564 96 -2548
rect -50 -2641 -34 -2607
rect 34 -2641 50 -2607
rect -230 -2745 -196 -2683
rect 196 -2745 230 -2683
rect -230 -2779 -134 -2745
rect 134 -2779 230 -2745
<< viali >>
rect -34 2607 34 2641
rect -96 2372 -62 2548
rect 62 2372 96 2548
rect -34 2279 34 2313
rect -96 2044 -62 2220
rect 62 2044 96 2220
rect -34 1951 34 1985
rect -96 1716 -62 1892
rect 62 1716 96 1892
rect -34 1623 34 1657
rect -96 1388 -62 1564
rect 62 1388 96 1564
rect -34 1295 34 1329
rect -96 1060 -62 1236
rect 62 1060 96 1236
rect -34 967 34 1001
rect -96 732 -62 908
rect 62 732 96 908
rect -34 639 34 673
rect -96 404 -62 580
rect 62 404 96 580
rect -34 311 34 345
rect -96 76 -62 252
rect 62 76 96 252
rect -34 -17 34 17
rect -96 -252 -62 -76
rect 62 -252 96 -76
rect -34 -345 34 -311
rect -96 -580 -62 -404
rect 62 -580 96 -404
rect -34 -673 34 -639
rect -96 -908 -62 -732
rect 62 -908 96 -732
rect -34 -1001 34 -967
rect -96 -1236 -62 -1060
rect 62 -1236 96 -1060
rect -34 -1329 34 -1295
rect -96 -1564 -62 -1388
rect 62 -1564 96 -1388
rect -34 -1657 34 -1623
rect -96 -1892 -62 -1716
rect 62 -1892 96 -1716
rect -34 -1985 34 -1951
rect -96 -2220 -62 -2044
rect 62 -2220 96 -2044
rect -34 -2313 34 -2279
rect -96 -2548 -62 -2372
rect 62 -2548 96 -2372
rect -34 -2641 34 -2607
<< metal1 >>
rect -46 2641 46 2647
rect -46 2607 -34 2641
rect 34 2607 46 2641
rect -46 2601 46 2607
rect -102 2548 -56 2560
rect -102 2372 -96 2548
rect -62 2372 -56 2548
rect -102 2360 -56 2372
rect 56 2548 102 2560
rect 56 2372 62 2548
rect 96 2372 102 2548
rect 56 2360 102 2372
rect -46 2313 46 2319
rect -46 2279 -34 2313
rect 34 2279 46 2313
rect -46 2273 46 2279
rect -102 2220 -56 2232
rect -102 2044 -96 2220
rect -62 2044 -56 2220
rect -102 2032 -56 2044
rect 56 2220 102 2232
rect 56 2044 62 2220
rect 96 2044 102 2220
rect 56 2032 102 2044
rect -46 1985 46 1991
rect -46 1951 -34 1985
rect 34 1951 46 1985
rect -46 1945 46 1951
rect -102 1892 -56 1904
rect -102 1716 -96 1892
rect -62 1716 -56 1892
rect -102 1704 -56 1716
rect 56 1892 102 1904
rect 56 1716 62 1892
rect 96 1716 102 1892
rect 56 1704 102 1716
rect -46 1657 46 1663
rect -46 1623 -34 1657
rect 34 1623 46 1657
rect -46 1617 46 1623
rect -102 1564 -56 1576
rect -102 1388 -96 1564
rect -62 1388 -56 1564
rect -102 1376 -56 1388
rect 56 1564 102 1576
rect 56 1388 62 1564
rect 96 1388 102 1564
rect 56 1376 102 1388
rect -46 1329 46 1335
rect -46 1295 -34 1329
rect 34 1295 46 1329
rect -46 1289 46 1295
rect -102 1236 -56 1248
rect -102 1060 -96 1236
rect -62 1060 -56 1236
rect -102 1048 -56 1060
rect 56 1236 102 1248
rect 56 1060 62 1236
rect 96 1060 102 1236
rect 56 1048 102 1060
rect -46 1001 46 1007
rect -46 967 -34 1001
rect 34 967 46 1001
rect -46 961 46 967
rect -102 908 -56 920
rect -102 732 -96 908
rect -62 732 -56 908
rect -102 720 -56 732
rect 56 908 102 920
rect 56 732 62 908
rect 96 732 102 908
rect 56 720 102 732
rect -46 673 46 679
rect -46 639 -34 673
rect 34 639 46 673
rect -46 633 46 639
rect -102 580 -56 592
rect -102 404 -96 580
rect -62 404 -56 580
rect -102 392 -56 404
rect 56 580 102 592
rect 56 404 62 580
rect 96 404 102 580
rect 56 392 102 404
rect -46 345 46 351
rect -46 311 -34 345
rect 34 311 46 345
rect -46 305 46 311
rect -102 252 -56 264
rect -102 76 -96 252
rect -62 76 -56 252
rect -102 64 -56 76
rect 56 252 102 264
rect 56 76 62 252
rect 96 76 102 252
rect 56 64 102 76
rect -46 17 46 23
rect -46 -17 -34 17
rect 34 -17 46 17
rect -46 -23 46 -17
rect -102 -76 -56 -64
rect -102 -252 -96 -76
rect -62 -252 -56 -76
rect -102 -264 -56 -252
rect 56 -76 102 -64
rect 56 -252 62 -76
rect 96 -252 102 -76
rect 56 -264 102 -252
rect -46 -311 46 -305
rect -46 -345 -34 -311
rect 34 -345 46 -311
rect -46 -351 46 -345
rect -102 -404 -56 -392
rect -102 -580 -96 -404
rect -62 -580 -56 -404
rect -102 -592 -56 -580
rect 56 -404 102 -392
rect 56 -580 62 -404
rect 96 -580 102 -404
rect 56 -592 102 -580
rect -46 -639 46 -633
rect -46 -673 -34 -639
rect 34 -673 46 -639
rect -46 -679 46 -673
rect -102 -732 -56 -720
rect -102 -908 -96 -732
rect -62 -908 -56 -732
rect -102 -920 -56 -908
rect 56 -732 102 -720
rect 56 -908 62 -732
rect 96 -908 102 -732
rect 56 -920 102 -908
rect -46 -967 46 -961
rect -46 -1001 -34 -967
rect 34 -1001 46 -967
rect -46 -1007 46 -1001
rect -102 -1060 -56 -1048
rect -102 -1236 -96 -1060
rect -62 -1236 -56 -1060
rect -102 -1248 -56 -1236
rect 56 -1060 102 -1048
rect 56 -1236 62 -1060
rect 96 -1236 102 -1060
rect 56 -1248 102 -1236
rect -46 -1295 46 -1289
rect -46 -1329 -34 -1295
rect 34 -1329 46 -1295
rect -46 -1335 46 -1329
rect -102 -1388 -56 -1376
rect -102 -1564 -96 -1388
rect -62 -1564 -56 -1388
rect -102 -1576 -56 -1564
rect 56 -1388 102 -1376
rect 56 -1564 62 -1388
rect 96 -1564 102 -1388
rect 56 -1576 102 -1564
rect -46 -1623 46 -1617
rect -46 -1657 -34 -1623
rect 34 -1657 46 -1623
rect -46 -1663 46 -1657
rect -102 -1716 -56 -1704
rect -102 -1892 -96 -1716
rect -62 -1892 -56 -1716
rect -102 -1904 -56 -1892
rect 56 -1716 102 -1704
rect 56 -1892 62 -1716
rect 96 -1892 102 -1716
rect 56 -1904 102 -1892
rect -46 -1951 46 -1945
rect -46 -1985 -34 -1951
rect 34 -1985 46 -1951
rect -46 -1991 46 -1985
rect -102 -2044 -56 -2032
rect -102 -2220 -96 -2044
rect -62 -2220 -56 -2044
rect -102 -2232 -56 -2220
rect 56 -2044 102 -2032
rect 56 -2220 62 -2044
rect 96 -2220 102 -2044
rect 56 -2232 102 -2220
rect -46 -2279 46 -2273
rect -46 -2313 -34 -2279
rect 34 -2313 46 -2279
rect -46 -2319 46 -2313
rect -102 -2372 -56 -2360
rect -102 -2548 -96 -2372
rect -62 -2548 -56 -2372
rect -102 -2560 -56 -2548
rect 56 -2372 102 -2360
rect 56 -2548 62 -2372
rect 96 -2548 102 -2372
rect 56 -2560 102 -2548
rect -46 -2607 46 -2601
rect -46 -2641 -34 -2607
rect 34 -2641 46 -2607
rect -46 -2647 46 -2641
<< properties >>
string FIXED_BBOX -213 -2762 213 2762
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.50 m 16 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
