magic
tech sky130A
timestamp 1666532281
<< metal4 >>
rect -154 4100 6 4101
rect -2956 1400 2956 4100
rect -2956 -1350 2956 1350
rect -2956 -4100 2956 -1400
rect -156 -4103 10 -4100
<< mimcap2 >>
rect -2906 4030 -306 4050
rect -2906 1470 -2886 4030
rect -326 1470 -306 4030
rect -2906 1450 -306 1470
rect 55 4030 2655 4050
rect 55 1470 75 4030
rect 2635 1470 2655 4030
rect 55 1450 2655 1470
rect -2906 1280 -306 1300
rect -2906 -1280 -2886 1280
rect -326 -1280 -306 1280
rect -2906 -1300 -306 -1280
rect 55 1280 2655 1300
rect 55 -1280 75 1280
rect 2635 -1280 2655 1280
rect 55 -1300 2655 -1280
rect -2906 -1470 -306 -1450
rect -2906 -4030 -2886 -1470
rect -326 -4030 -306 -1470
rect -2906 -4050 -306 -4030
rect 55 -1470 2655 -1450
rect 55 -4030 75 -1470
rect 2635 -4030 2655 -1470
rect 55 -4050 2655 -4030
<< mimcap2contact >>
rect -2886 1470 -326 4030
rect 75 1470 2635 4030
rect -2886 -1280 -326 1280
rect 75 -1280 2635 1280
rect -2886 -4030 -326 -1470
rect 75 -4030 2635 -1470
<< metal5 >>
rect -1686 4042 -1526 4125
rect -326 4042 -166 4125
rect 1275 4042 1435 4125
rect 2635 4042 2795 4125
rect -2898 4030 -166 4042
rect -2898 1470 -2886 4030
rect -326 1470 -166 4030
rect -2898 1458 -166 1470
rect 63 4030 2795 4042
rect 63 1470 75 4030
rect 2635 1470 2795 4030
rect 63 1458 2795 1470
rect -1686 1292 -1526 1458
rect -326 1292 -166 1458
rect 1275 1292 1435 1458
rect 2635 1292 2795 1458
rect -2898 1280 -166 1292
rect -2898 -1280 -2886 1280
rect -326 -1280 -166 1280
rect -2898 -1292 -166 -1280
rect 63 1280 2795 1292
rect 63 -1280 75 1280
rect 2635 -1280 2795 1280
rect 63 -1292 2795 -1280
rect -1686 -1458 -1526 -1292
rect -326 -1458 -166 -1292
rect 1275 -1458 1435 -1292
rect 2635 -1458 2795 -1292
rect -2898 -1470 -166 -1458
rect -2898 -4030 -2886 -1470
rect -326 -4030 -166 -1470
rect -2898 -4042 -166 -4030
rect 63 -1470 2795 -1458
rect 63 -4030 75 -1470
rect 2635 -4030 2795 -1470
rect 63 -4042 2795 -4030
rect -1686 -4125 -1526 -4042
rect -326 -4125 -166 -4042
rect 1275 -4125 1435 -4042
rect 2635 -4125 2795 -4042
<< properties >>
string FIXED_BBOX 5 1400 2705 4100
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 26.00 l 26.00 val 1.371k carea 2.00 cperi 0.19 nx 2 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
