magic
tech sky130A
magscale 1 2
timestamp 1666205007
<< nwell >>
rect -246 -4219 246 4219
<< pmos >>
rect -50 -4000 50 4000
<< pdiff >>
rect -108 3988 -50 4000
rect -108 -3988 -96 3988
rect -62 -3988 -50 3988
rect -108 -4000 -50 -3988
rect 50 3988 108 4000
rect 50 -3988 62 3988
rect 96 -3988 108 3988
rect 50 -4000 108 -3988
<< pdiffc >>
rect -96 -3988 -62 3988
rect 62 -3988 96 3988
<< nsubdiff >>
rect -210 4149 -114 4183
rect 114 4149 210 4183
rect -210 4087 -176 4149
rect 176 4087 210 4149
rect -210 -4149 -176 -4087
rect 176 -4149 210 -4087
rect -210 -4183 -114 -4149
rect 114 -4183 210 -4149
<< nsubdiffcont >>
rect -114 4149 114 4183
rect -210 -4087 -176 4087
rect 176 -4087 210 4087
rect -114 -4183 114 -4149
<< poly >>
rect -50 4081 50 4097
rect -50 4047 -34 4081
rect 34 4047 50 4081
rect -50 4000 50 4047
rect -50 -4047 50 -4000
rect -50 -4081 -34 -4047
rect 34 -4081 50 -4047
rect -50 -4097 50 -4081
<< polycont >>
rect -34 4047 34 4081
rect -34 -4081 34 -4047
<< locali >>
rect -210 4149 -114 4183
rect 114 4149 210 4183
rect -210 4087 -176 4149
rect 176 4087 210 4149
rect -50 4047 -34 4081
rect 34 4047 50 4081
rect -96 3988 -62 4004
rect -96 -4004 -62 -3988
rect 62 3988 96 4004
rect 62 -4004 96 -3988
rect -50 -4081 -34 -4047
rect 34 -4081 50 -4047
rect -210 -4149 -176 -4087
rect 176 -4149 210 -4087
rect -210 -4183 -114 -4149
rect 114 -4183 210 -4149
<< viali >>
rect -34 4047 34 4081
rect -96 -3988 -62 3988
rect 62 -3988 96 3988
rect -34 -4081 34 -4047
<< metal1 >>
rect -46 4081 46 4087
rect -46 4047 -34 4081
rect 34 4047 46 4081
rect -46 4041 46 4047
rect -102 3988 -56 4000
rect -102 -3988 -96 3988
rect -62 -3988 -56 3988
rect -102 -4000 -56 -3988
rect 56 3988 102 4000
rect 56 -3988 62 3988
rect 96 -3988 102 3988
rect 56 -4000 102 -3988
rect -46 -4047 46 -4041
rect -46 -4081 -34 -4047
rect 34 -4081 46 -4047
rect -46 -4087 46 -4081
<< properties >>
string FIXED_BBOX -193 -4166 193 4166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 40 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
