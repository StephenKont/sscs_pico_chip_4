magic
tech sky130A
magscale 1 2
timestamp 1668298669
<< viali >>
rect 15407 17976 18271 18010
rect 15311 6674 15345 17914
rect 15617 17766 16665 17800
rect 17013 17766 18061 17800
rect 15521 16656 15555 17704
rect 16727 16656 16761 17704
rect 16917 16656 16951 17704
rect 18123 16656 18157 17704
rect 15617 16560 16665 16594
rect 17013 16560 18061 16594
rect 15617 16370 16665 16404
rect 17013 16370 18061 16404
rect 15521 15260 15555 16308
rect 16727 15260 16761 16308
rect 16917 15260 16951 16308
rect 18123 15260 18157 16308
rect 15617 15164 16665 15198
rect 17013 15164 18061 15198
rect 15617 14974 16665 15008
rect 17013 14974 18061 15008
rect 15521 13864 15555 14912
rect 16727 13864 16761 14912
rect 16917 13864 16951 14912
rect 18123 13864 18157 14912
rect 15617 13768 16665 13802
rect 17013 13768 18061 13802
rect 15617 13578 16665 13612
rect 17013 13578 18061 13612
rect 15521 12468 15555 13516
rect 16727 12468 16761 13516
rect 16917 12468 16951 13516
rect 18123 12468 18157 13516
rect 15617 12372 16665 12406
rect 17013 12372 18061 12406
rect 15617 12182 16665 12216
rect 17013 12182 18061 12216
rect 15521 11072 15555 12120
rect 16727 11072 16761 12120
rect 16917 11072 16951 12120
rect 18123 11072 18157 12120
rect 15617 10976 16665 11010
rect 17013 10976 18061 11010
rect 15617 10786 16665 10820
rect 17013 10786 18061 10820
rect 15521 9676 15555 10724
rect 16727 9676 16761 10724
rect 16917 9676 16951 10724
rect 18123 9676 18157 10724
rect 15617 9580 16665 9614
rect 17013 9580 18061 9614
rect 15617 9390 16665 9424
rect 17013 9390 18061 9424
rect 15521 8280 15555 9328
rect 16727 8280 16761 9328
rect 16917 8280 16951 9328
rect 18123 8280 18157 9328
rect 15617 8184 16665 8218
rect 17013 8184 18061 8218
rect 15617 7994 16665 8028
rect 17013 7994 18061 8028
rect 15521 6884 15555 7932
rect 16727 6884 16761 7932
rect 16917 6884 16951 7932
rect 18123 6884 18157 7932
rect 15617 6788 16665 6822
rect 17013 6788 18061 6822
rect 18333 6674 18367 17914
rect 15407 6578 18271 6612
rect 5116 5038 6198 5072
rect 6260 4838 6294 4976
rect 5624 4742 6198 4776
rect 15388 2373 16542 2407
rect 15292 2173 15326 2311
rect 16604 2173 16638 2311
rect 15388 2077 16542 2111
rect 15388 1655 16542 1689
rect 15292 1455 15326 1593
rect 16604 1455 16638 1593
rect 15388 1359 16542 1393
rect 8712 982 9888 1016
rect 10154 966 11236 1000
rect 8616 570 8650 920
rect 9950 570 9984 920
rect 10058 766 10092 904
rect 11298 766 11332 904
rect 10154 670 11236 704
rect 8712 474 9888 508
<< metal1 >>
rect 16714 19074 16964 19086
rect 16714 18811 16726 19074
rect 16952 18811 16964 19074
rect 16714 18022 16964 18811
rect 15299 18010 18379 18022
rect 15299 17976 15407 18010
rect 18271 17976 18379 18010
rect 15299 17964 18379 17976
rect 15299 17914 15357 17964
rect 15299 6674 15311 17914
rect 15345 6674 15357 17914
rect 18321 17914 18379 17964
rect 15443 17800 18235 17878
rect 15443 17766 15617 17800
rect 16665 17766 17013 17800
rect 18061 17766 18235 17800
rect 15443 17754 18235 17766
rect 15443 17704 15567 17754
rect 15443 16656 15521 17704
rect 15555 16656 15567 17704
rect 16715 17704 16963 17754
rect 15443 16606 15567 16656
rect 16715 16656 16727 17704
rect 16761 16656 16917 17704
rect 16951 16656 16963 17704
rect 18111 17704 18235 17754
rect 16715 16606 16963 16656
rect 18111 16656 18123 17704
rect 18157 16656 18235 17704
rect 18111 16606 18235 16656
rect 15443 16596 18235 16606
rect 15443 16368 15453 16596
rect 18221 16368 18235 16596
rect 15443 16358 18235 16368
rect 15443 16308 15567 16358
rect 15443 15260 15521 16308
rect 15555 15260 15567 16308
rect 16715 16308 16963 16358
rect 15443 15210 15567 15260
rect 16715 15260 16727 16308
rect 16761 15260 16917 16308
rect 16951 15260 16963 16308
rect 18111 16308 18235 16358
rect 16715 15210 16963 15260
rect 18111 15260 18123 16308
rect 18157 15260 18235 16308
rect 18111 15210 18235 15260
rect 15443 15200 18235 15210
rect 15443 14972 15453 15200
rect 18221 14972 18235 15200
rect 15443 14962 18235 14972
rect 15443 14912 15567 14962
rect 15443 13864 15521 14912
rect 15555 13864 15567 14912
rect 16715 14912 16963 14962
rect 15443 13814 15567 13864
rect 16715 13864 16727 14912
rect 16761 13864 16917 14912
rect 16951 13864 16963 14912
rect 18111 14912 18235 14962
rect 16715 13814 16963 13864
rect 18111 13864 18123 14912
rect 18157 13864 18235 14912
rect 18111 13814 18235 13864
rect 15443 13804 18235 13814
rect 15443 13576 15453 13804
rect 18221 13576 18235 13804
rect 15443 13566 18235 13576
rect 15443 13516 15567 13566
rect 15443 12468 15521 13516
rect 15555 12468 15567 13516
rect 16715 13516 16963 13566
rect 15443 12418 15567 12468
rect 16715 12468 16727 13516
rect 16761 12468 16917 13516
rect 16951 12468 16963 13516
rect 18111 13516 18235 13566
rect 16715 12418 16963 12468
rect 18111 12468 18123 13516
rect 18157 12468 18235 13516
rect 18111 12418 18235 12468
rect 15443 12408 18235 12418
rect 15443 12180 15453 12408
rect 18221 12180 18235 12408
rect 15443 12170 18235 12180
rect 15443 12120 15567 12170
rect 15443 11072 15521 12120
rect 15555 11072 15567 12120
rect 16715 12120 16963 12170
rect 15443 11022 15567 11072
rect 16715 11072 16727 12120
rect 16761 11072 16917 12120
rect 16951 11072 16963 12120
rect 18111 12120 18235 12170
rect 16715 11022 16963 11072
rect 18111 11072 18123 12120
rect 18157 11072 18235 12120
rect 18111 11022 18235 11072
rect 15443 11012 18235 11022
rect 15443 10784 15453 11012
rect 18221 10784 18235 11012
rect 15443 10774 18235 10784
rect 15443 10724 15567 10774
rect 15443 9676 15521 10724
rect 15555 9676 15567 10724
rect 16715 10724 16963 10774
rect 15443 9626 15567 9676
rect 16715 9676 16727 10724
rect 16761 9676 16917 10724
rect 16951 9676 16963 10724
rect 18111 10724 18235 10774
rect 16715 9626 16963 9676
rect 18111 9676 18123 10724
rect 18157 9676 18235 10724
rect 18111 9626 18235 9676
rect 15443 9616 18235 9626
rect 15443 9388 15453 9616
rect 18221 9388 18235 9616
rect 15443 9378 18235 9388
rect 15443 9328 15567 9378
rect 15443 8280 15521 9328
rect 15555 8280 15567 9328
rect 16715 9328 16963 9378
rect 15443 8230 15567 8280
rect 16715 8280 16727 9328
rect 16761 8280 16917 9328
rect 16951 8280 16963 9328
rect 18111 9328 18235 9378
rect 16715 8230 16963 8280
rect 18111 8280 18123 9328
rect 18157 8280 18235 9328
rect 18111 8230 18235 8280
rect 15443 8220 18235 8230
rect 15443 7992 15453 8220
rect 18221 7992 18235 8220
rect 15443 7982 18235 7992
rect 15443 7932 15567 7982
rect 15443 6884 15521 7932
rect 15555 6884 15567 7932
rect 16715 7932 16963 7982
rect 15443 6834 15567 6884
rect 16715 6884 16727 7932
rect 16761 6884 16917 7932
rect 16951 6884 16963 7932
rect 18111 7932 18235 7982
rect 16715 6834 16963 6884
rect 18111 6884 18123 7932
rect 18157 6884 18235 7932
rect 18111 6834 18235 6884
rect 15443 6822 18235 6834
rect 15443 6788 15617 6822
rect 16665 6788 17013 6822
rect 18061 6788 18235 6822
rect 15443 6710 18235 6788
rect 15299 6624 15357 6674
rect 18321 6674 18333 17914
rect 18367 6674 18379 17914
rect 18321 6624 18379 6674
rect 15299 6612 18379 6624
rect 15299 6578 15407 6612
rect 18271 6578 18379 6612
rect 15299 6566 18379 6578
rect 16716 6530 16964 6566
rect 7098 5527 12654 5552
rect 7098 5334 7124 5527
rect 12624 5334 12654 5527
rect 7098 5310 12654 5334
rect 5020 5072 6301 5080
rect 5020 5038 5116 5072
rect 6198 5038 6301 5072
rect 5020 5031 6301 5038
rect 6253 4976 6301 5031
rect 4502 4742 5582 4942
rect 5732 4936 6164 4942
rect 5732 4878 5738 4936
rect 6158 4878 6164 4936
rect 5732 4872 6164 4878
rect 6253 4838 6260 4976
rect 6294 4838 6301 4976
rect 6253 4789 6301 4838
rect 5612 4776 6301 4789
rect 5612 4742 5624 4776
rect 6198 4742 6301 4776
rect 4502 2580 4702 4742
rect 5612 4730 6301 4742
rect 5616 4624 5737 4730
rect 5616 4527 5622 4624
rect 5731 4527 5737 4624
rect 5616 4522 5737 4527
rect 6722 4629 9772 4719
rect 4876 4143 5012 4151
rect 4876 4050 4885 4143
rect 5003 4133 5012 4143
rect 6722 4133 6812 4629
rect 5003 4050 6812 4133
rect 4876 4043 6812 4050
rect 4876 4042 4974 4043
rect 4502 2298 4508 2580
rect 4692 2382 4702 2580
rect 9682 2382 9772 4629
rect 15255 2407 16662 2431
rect 4692 2298 4918 2382
rect 4502 2292 4918 2298
rect 9682 2292 9950 2382
rect 15255 2373 15388 2407
rect 16542 2373 16662 2407
rect 15255 2358 16662 2373
rect 15255 2311 15339 2358
rect 9632 2242 9954 2248
rect 9632 2162 9638 2242
rect 9786 2162 9954 2242
rect 9632 2156 9954 2162
rect 15255 2173 15292 2311
rect 15326 2173 15339 2311
rect 16583 2311 16662 2358
rect 15422 2270 15854 2277
rect 15422 2214 15429 2270
rect 15846 2214 15854 2270
rect 15422 2207 15854 2214
rect 16076 2270 16508 2278
rect 16076 2218 16084 2270
rect 16498 2218 16508 2270
rect 16076 2208 16508 2218
rect 15255 2130 15339 2173
rect 16583 2173 16604 2311
rect 16638 2173 16662 2311
rect 16583 2130 16662 2173
rect 15255 2111 16662 2130
rect 15255 2077 15388 2111
rect 16542 2077 16662 2111
rect 15255 2053 16662 2077
rect 15255 1713 15339 2053
rect 16392 1713 16450 2053
rect 15255 1689 16662 1713
rect 15255 1655 15388 1689
rect 16542 1655 16662 1689
rect 4751 1630 4835 1640
rect 4751 1561 4760 1630
rect 4825 1618 4835 1630
rect 15255 1635 16662 1655
rect 4825 1561 4982 1618
rect 4751 1554 4982 1561
rect 7094 1390 7554 1615
rect 11296 1590 12628 1616
rect 6393 1345 7554 1390
rect 6393 724 6452 1345
rect 7488 724 7554 1345
rect 10394 1546 12628 1590
rect 10394 1164 10460 1546
rect 11242 1390 12628 1546
rect 15255 1593 15339 1635
rect 15255 1455 15292 1593
rect 15326 1455 15339 1593
rect 16589 1593 16662 1635
rect 15422 1551 15854 1559
rect 15422 1496 15430 1551
rect 15845 1496 15854 1551
rect 15422 1489 15854 1496
rect 15255 1414 15339 1455
rect 16076 1414 16508 1559
rect 16589 1455 16604 1593
rect 16638 1455 16662 1593
rect 16589 1414 16662 1455
rect 15255 1393 16662 1414
rect 11242 1164 11301 1390
rect 10394 1119 11301 1164
rect 6393 680 7554 724
rect 8580 1036 10020 1052
rect 12160 1036 12240 1390
rect 12534 1282 12618 1390
rect 15255 1359 15388 1393
rect 16542 1359 16662 1393
rect 15255 1335 16662 1359
rect 15255 1282 15339 1335
rect 12534 1198 15339 1282
rect 8580 1016 12240 1036
rect 8580 982 8712 1016
rect 9888 1000 12240 1016
rect 9888 982 10154 1000
rect 8580 972 10154 982
rect 8580 920 8660 972
rect 8580 570 8616 920
rect 8650 570 8660 920
rect 9940 966 10154 972
rect 11236 966 12240 1000
rect 9940 956 12240 966
rect 9940 920 10103 956
rect 8580 518 8660 570
rect 9940 570 9950 920
rect 9984 904 10103 920
rect 9984 766 10058 904
rect 10092 766 10103 904
rect 11285 904 11368 956
rect 10188 864 10620 870
rect 10188 806 10194 864
rect 10614 806 10620 864
rect 10188 800 10620 806
rect 10770 864 11202 870
rect 10770 806 10776 864
rect 11196 806 11202 864
rect 10770 800 11202 806
rect 9984 714 10103 766
rect 11285 766 11298 904
rect 11332 766 11368 904
rect 11285 714 11368 766
rect 9984 704 11368 714
rect 9984 670 10154 704
rect 11236 670 11368 704
rect 9984 634 11368 670
rect 9984 570 10020 634
rect 9940 518 10020 570
rect 8580 508 10020 518
rect 8580 474 8712 508
rect 9888 474 10020 508
rect 8580 438 10020 474
rect 11406 -326 11591 -316
rect 11406 -491 11416 -326
rect 11580 -491 11591 -326
rect 11406 -501 11591 -491
rect 11498 -1220 11591 -501
rect 11498 -1312 11647 -1220
rect 13704 -2051 14611 -2007
rect 13704 -2433 13770 -2051
rect 14552 -2433 14611 -2051
rect 13704 -2478 14611 -2433
<< via1 >>
rect 16726 18811 16952 19074
rect 15841 16880 16441 17480
rect 17237 16880 17837 17480
rect 15453 16594 18221 16596
rect 15453 16560 15617 16594
rect 15617 16560 16665 16594
rect 16665 16560 17013 16594
rect 17013 16560 18061 16594
rect 18061 16560 18221 16594
rect 15453 16404 18221 16560
rect 15453 16370 15617 16404
rect 15617 16370 16665 16404
rect 16665 16370 17013 16404
rect 17013 16370 18061 16404
rect 18061 16370 18221 16404
rect 15453 16368 18221 16370
rect 15841 15484 16441 16084
rect 17237 15484 17837 16084
rect 15453 15198 18221 15200
rect 15453 15164 15617 15198
rect 15617 15164 16665 15198
rect 16665 15164 17013 15198
rect 17013 15164 18061 15198
rect 18061 15164 18221 15198
rect 15453 15008 18221 15164
rect 15453 14974 15617 15008
rect 15617 14974 16665 15008
rect 16665 14974 17013 15008
rect 17013 14974 18061 15008
rect 18061 14974 18221 15008
rect 15453 14972 18221 14974
rect 15841 14088 16441 14688
rect 17237 14088 17837 14688
rect 15453 13802 18221 13804
rect 15453 13768 15617 13802
rect 15617 13768 16665 13802
rect 16665 13768 17013 13802
rect 17013 13768 18061 13802
rect 18061 13768 18221 13802
rect 15453 13612 18221 13768
rect 15453 13578 15617 13612
rect 15617 13578 16665 13612
rect 16665 13578 17013 13612
rect 17013 13578 18061 13612
rect 18061 13578 18221 13612
rect 15453 13576 18221 13578
rect 15841 12692 16441 13292
rect 17237 12692 17837 13292
rect 15453 12406 18221 12408
rect 15453 12372 15617 12406
rect 15617 12372 16665 12406
rect 16665 12372 17013 12406
rect 17013 12372 18061 12406
rect 18061 12372 18221 12406
rect 15453 12216 18221 12372
rect 15453 12182 15617 12216
rect 15617 12182 16665 12216
rect 16665 12182 17013 12216
rect 17013 12182 18061 12216
rect 18061 12182 18221 12216
rect 15453 12180 18221 12182
rect 15841 11296 16441 11896
rect 17237 11296 17837 11896
rect 15453 11010 18221 11012
rect 15453 10976 15617 11010
rect 15617 10976 16665 11010
rect 16665 10976 17013 11010
rect 17013 10976 18061 11010
rect 18061 10976 18221 11010
rect 15453 10820 18221 10976
rect 15453 10786 15617 10820
rect 15617 10786 16665 10820
rect 16665 10786 17013 10820
rect 17013 10786 18061 10820
rect 18061 10786 18221 10820
rect 15453 10784 18221 10786
rect 15841 9900 16441 10500
rect 17237 9900 17837 10500
rect 15453 9614 18221 9616
rect 15453 9580 15617 9614
rect 15617 9580 16665 9614
rect 16665 9580 17013 9614
rect 17013 9580 18061 9614
rect 18061 9580 18221 9614
rect 15453 9424 18221 9580
rect 15453 9390 15617 9424
rect 15617 9390 16665 9424
rect 16665 9390 17013 9424
rect 17013 9390 18061 9424
rect 18061 9390 18221 9424
rect 15453 9388 18221 9390
rect 15841 8504 16441 9104
rect 17237 8504 17837 9104
rect 15453 8218 18221 8220
rect 15453 8184 15617 8218
rect 15617 8184 16665 8218
rect 16665 8184 17013 8218
rect 17013 8184 18061 8218
rect 18061 8184 18221 8218
rect 15453 8028 18221 8184
rect 15453 7994 15617 8028
rect 15617 7994 16665 8028
rect 16665 7994 17013 8028
rect 17013 7994 18061 8028
rect 18061 7994 18221 8028
rect 15453 7992 18221 7994
rect 15841 7108 16441 7708
rect 17237 7108 17837 7708
rect 7124 5334 12624 5527
rect 5738 4878 6158 4936
rect 5622 4527 5731 4624
rect 4885 4050 5003 4143
rect 4508 2298 4692 2580
rect 4885 2166 4964 2239
rect 9638 2162 9786 2242
rect 15429 2214 15846 2270
rect 16084 2218 16498 2270
rect 4760 1561 4825 1630
rect 6452 724 7488 1345
rect 10460 1164 11242 1546
rect 15430 1496 15845 1551
rect 8758 620 9010 864
rect 9440 620 9836 870
rect 10194 806 10614 864
rect 10776 806 11196 864
rect 11416 -491 11580 -326
rect 13770 -2433 14552 -2051
<< metal2 >>
rect 4555 19074 16964 19086
rect 4555 19057 16726 19074
rect 4555 5954 4575 19057
rect 4814 18811 16726 19057
rect 16952 18811 16964 19074
rect 4814 18801 16964 18811
rect 4814 18314 4840 18801
rect 14929 18472 15258 18480
rect 14832 18450 15258 18472
rect 14832 18424 14963 18450
rect 4814 18266 4920 18314
rect 4814 17998 4840 18266
rect 14929 18156 14963 18424
rect 14832 18108 14963 18156
rect 4814 17950 4920 17998
rect 4814 17682 4840 17950
rect 14929 17840 14963 18108
rect 14832 17792 14963 17840
rect 4814 17634 4920 17682
rect 4814 17366 4840 17634
rect 14929 17524 14963 17792
rect 14832 17476 14963 17524
rect 4814 17318 4920 17366
rect 4814 17050 4840 17318
rect 14929 17208 14963 17476
rect 14832 17160 14963 17208
rect 4814 17002 4920 17050
rect 4814 16734 4840 17002
rect 14929 16892 14963 17160
rect 14832 16844 14963 16892
rect 4814 16686 4920 16734
rect 4814 16418 4840 16686
rect 14929 16576 14963 16844
rect 14832 16528 14963 16576
rect 4814 16370 4920 16418
rect 4814 16102 4840 16370
rect 14929 16260 14963 16528
rect 14832 16212 14963 16260
rect 4814 16054 4920 16102
rect 4814 15786 4840 16054
rect 14929 15944 14963 16212
rect 14832 15896 14963 15944
rect 4814 15738 4920 15786
rect 4814 15470 4840 15738
rect 14929 15628 14963 15896
rect 14832 15580 14963 15628
rect 4814 15422 4920 15470
rect 4814 15154 4840 15422
rect 14929 15312 14963 15580
rect 14832 15264 14963 15312
rect 4814 15106 4920 15154
rect 4814 14838 4840 15106
rect 14929 14996 14963 15264
rect 14832 14948 14963 14996
rect 4814 14790 4920 14838
rect 4814 14522 4840 14790
rect 14929 14680 14963 14948
rect 14832 14632 14963 14680
rect 4814 14474 4920 14522
rect 4814 14206 4840 14474
rect 14929 14364 14963 14632
rect 14832 14316 14963 14364
rect 4814 14158 4920 14206
rect 4814 13890 4840 14158
rect 14929 14048 14963 14316
rect 14832 14000 14963 14048
rect 4814 13842 4920 13890
rect 4814 13574 4840 13842
rect 14929 13732 14963 14000
rect 14832 13684 14963 13732
rect 4814 13526 4920 13574
rect 4814 13258 4840 13526
rect 14929 13416 14963 13684
rect 14832 13368 14963 13416
rect 4814 13210 4920 13258
rect 4814 12942 4840 13210
rect 14929 13100 14963 13368
rect 14832 13052 14963 13100
rect 4814 12894 4920 12942
rect 4814 12626 4840 12894
rect 14929 12784 14963 13052
rect 14832 12736 14963 12784
rect 4814 12578 4920 12626
rect 4814 12310 4840 12578
rect 14929 12468 14963 12736
rect 14832 12420 14963 12468
rect 4814 12262 4920 12310
rect 4814 11994 4840 12262
rect 14929 12152 14963 12420
rect 14832 12104 14963 12152
rect 4814 11946 4920 11994
rect 4814 11678 4840 11946
rect 14929 11836 14963 12104
rect 14832 11788 14963 11836
rect 4814 11630 4920 11678
rect 4814 11362 4840 11630
rect 14929 11520 14963 11788
rect 14832 11472 14963 11520
rect 4814 11314 4920 11362
rect 4814 11046 4840 11314
rect 14929 11204 14963 11472
rect 14832 11156 14963 11204
rect 4814 10998 4920 11046
rect 4814 10730 4840 10998
rect 14929 10888 14963 11156
rect 14832 10840 14963 10888
rect 4814 10682 4920 10730
rect 4814 10414 4840 10682
rect 14929 10572 14963 10840
rect 14832 10524 14963 10572
rect 4814 10366 4920 10414
rect 4814 10098 4840 10366
rect 14929 10256 14963 10524
rect 14832 10208 14963 10256
rect 4814 10050 4920 10098
rect 4814 9782 4840 10050
rect 14929 9940 14963 10208
rect 14832 9892 14963 9940
rect 4814 9734 4920 9782
rect 4814 9466 4840 9734
rect 14929 9624 14963 9892
rect 14832 9576 14963 9624
rect 4814 9418 4920 9466
rect 4814 9150 4840 9418
rect 14929 9308 14963 9576
rect 14832 9260 14963 9308
rect 4814 9102 4920 9150
rect 4814 8834 4840 9102
rect 14929 8992 14963 9260
rect 14832 8944 14963 8992
rect 4814 8786 4920 8834
rect 4814 8518 4840 8786
rect 14929 8676 14963 8944
rect 14832 8628 14963 8676
rect 4814 8470 4920 8518
rect 4814 8202 4840 8470
rect 14929 8360 14963 8628
rect 14832 8312 14963 8360
rect 4814 8154 4920 8202
rect 4814 7886 4840 8154
rect 14929 8044 14963 8312
rect 14832 7996 14963 8044
rect 4814 7838 4920 7886
rect 4814 7570 4840 7838
rect 14929 7728 14963 7996
rect 14832 7680 14963 7728
rect 4814 7522 4920 7570
rect 4814 7254 4840 7522
rect 14929 7412 14963 7680
rect 14832 7364 14963 7412
rect 4814 7206 4920 7254
rect 4814 6938 4840 7206
rect 14929 7096 14963 7364
rect 14832 7048 14963 7096
rect 4814 6890 4920 6938
rect 4814 6622 4840 6890
rect 14929 6780 14963 7048
rect 14832 6732 14963 6780
rect 4814 6574 4920 6622
rect 4814 6306 4840 6574
rect 14929 6464 14963 6732
rect 14832 6416 14963 6464
rect 4814 6258 4920 6306
rect 4814 5990 4840 6258
rect 14929 6148 14963 6416
rect 14832 6100 14963 6148
rect 4814 5954 4920 5990
rect 4555 5942 4920 5954
rect 4555 5933 4840 5942
rect 14929 5832 14963 6100
rect 14832 5804 14963 5832
rect 15226 17480 15258 18450
rect 15741 17480 16541 17580
rect 17137 17480 17937 17580
rect 15226 16880 15841 17480
rect 16441 16880 17237 17480
rect 17837 16880 17937 17480
rect 15226 16084 15258 16880
rect 15741 16780 16541 16880
rect 17137 16780 17937 16880
rect 15443 16596 18637 16606
rect 15443 16368 15453 16596
rect 18221 16368 18637 16596
rect 15443 16358 18637 16368
rect 15741 16084 16541 16184
rect 17137 16084 17937 16184
rect 15226 15484 15841 16084
rect 16441 15484 17237 16084
rect 17837 15484 17937 16084
rect 15226 14688 15258 15484
rect 15741 15384 16541 15484
rect 17137 15384 17937 15484
rect 18463 15210 18637 16358
rect 15443 15200 18637 15210
rect 15443 14972 15453 15200
rect 18221 14972 18637 15200
rect 15443 14962 18637 14972
rect 15741 14688 16541 14788
rect 17137 14688 17937 14788
rect 15226 14088 15841 14688
rect 16441 14088 17237 14688
rect 17837 14088 17937 14688
rect 15226 13292 15258 14088
rect 15741 13988 16541 14088
rect 17137 13988 17937 14088
rect 18463 13814 18637 14962
rect 15443 13804 18637 13814
rect 15443 13576 15453 13804
rect 18221 13576 18637 13804
rect 15443 13566 18637 13576
rect 15741 13292 16541 13392
rect 17137 13292 17937 13392
rect 15226 12692 15841 13292
rect 16441 12692 17237 13292
rect 17837 12692 17937 13292
rect 15226 11896 15258 12692
rect 15741 12592 16541 12692
rect 17137 12592 17937 12692
rect 18463 12418 18637 13566
rect 15443 12408 18637 12418
rect 15443 12180 15453 12408
rect 18221 12180 18637 12408
rect 15443 12170 18637 12180
rect 15741 11896 16541 11996
rect 17137 11896 17937 11996
rect 15226 11296 15841 11896
rect 16441 11296 17237 11896
rect 17837 11296 17937 11896
rect 15226 10500 15258 11296
rect 15741 11196 16541 11296
rect 17137 11196 17937 11296
rect 18463 11022 18637 12170
rect 15443 11012 18637 11022
rect 15443 10784 15453 11012
rect 18221 10784 18637 11012
rect 15443 10774 18637 10784
rect 15741 10500 16541 10600
rect 17137 10500 17937 10600
rect 15226 9900 15841 10500
rect 16441 9900 17237 10500
rect 17837 9900 17937 10500
rect 15226 9104 15258 9900
rect 15741 9800 16541 9900
rect 17137 9800 17937 9900
rect 18463 9626 18637 10774
rect 15443 9616 18637 9626
rect 15443 9388 15453 9616
rect 18221 9388 18637 9616
rect 15443 9378 18637 9388
rect 15741 9104 16541 9204
rect 17137 9104 17937 9204
rect 15226 8504 15841 9104
rect 16441 8504 17237 9104
rect 17837 8504 17937 9104
rect 15226 7708 15258 8504
rect 15741 8404 16541 8504
rect 17137 8404 17937 8504
rect 18463 8230 18637 9378
rect 15443 8220 18637 8230
rect 15443 7992 15453 8220
rect 18221 7992 18637 8220
rect 15443 7982 18637 7992
rect 15741 7708 16541 7808
rect 17137 7708 17937 7808
rect 15226 7108 15841 7708
rect 16441 7108 17237 7708
rect 17837 7108 17937 7708
rect 15226 5804 15258 7108
rect 15741 7008 16541 7108
rect 17137 7008 17937 7108
rect 18463 6128 18637 7982
rect 14832 5784 15258 5804
rect 14929 5776 15258 5784
rect 16452 5954 18637 6128
rect 7098 5527 12654 5552
rect 7098 5334 7124 5527
rect 12624 5334 12654 5527
rect 7098 5070 7152 5334
rect 12579 5070 12654 5334
rect 7098 5019 12654 5070
rect 5726 4936 6170 4948
rect 5726 4878 5738 4936
rect 6158 4878 6170 4936
rect 5726 4866 6170 4878
rect 14903 4820 15493 4824
rect 14340 4818 15498 4820
rect 8342 4815 15556 4818
rect 5616 4624 5737 4631
rect 5616 4606 5622 4624
rect 4751 4527 5622 4606
rect 5731 4527 5737 4624
rect 4751 4522 5737 4527
rect 4498 2580 4702 2588
rect 4498 2298 4508 2580
rect 4692 2298 4702 2580
rect 4498 2288 4702 2298
rect 4751 1630 4835 4522
rect 8342 4225 14903 4815
rect 15493 4225 15556 4815
rect 8342 4218 15556 4225
rect 4876 4143 5012 4151
rect 4876 4050 4885 4143
rect 5003 4050 5012 4143
rect 4876 4043 5012 4050
rect 4876 4042 4974 4043
rect 8342 3886 8942 4218
rect 13416 3952 14016 4218
rect 14903 4216 15493 4218
rect 16452 2838 16626 5954
rect 16240 2664 16626 2838
rect 16240 2278 16414 2664
rect 15422 2270 15854 2277
rect 4876 2239 4974 2248
rect 4876 2166 4885 2239
rect 4964 2166 4974 2239
rect 4876 2156 4974 2166
rect 9632 2242 9794 2248
rect 9632 2162 9638 2242
rect 9786 2162 9794 2242
rect 4751 1561 4760 1630
rect 4825 1561 4835 1630
rect 4751 1554 4835 1561
rect 9632 1944 9794 2162
rect 15422 2214 15429 2270
rect 15846 2214 15854 2270
rect 6393 1345 7554 1390
rect 6393 724 6452 1345
rect 7488 724 7554 1345
rect 6393 680 7554 724
rect 8752 864 9016 1442
rect 9632 876 9792 1944
rect 15422 1811 15854 2214
rect 16076 2270 16508 2278
rect 16076 2218 16084 2270
rect 16498 2218 16508 2270
rect 16076 2207 16508 2218
rect 15422 1626 15440 1811
rect 15836 1626 15854 1811
rect 10394 1546 11301 1590
rect 10394 1164 10460 1546
rect 11242 1536 11301 1546
rect 15422 1551 15854 1626
rect 11242 1390 12035 1536
rect 15422 1496 15430 1551
rect 15845 1496 15854 1551
rect 15422 1489 15854 1496
rect 11242 1164 11301 1390
rect 10394 1119 11301 1164
rect 13547 979 13617 1443
rect 11533 909 13617 979
rect 16122 999 16722 1034
rect 8752 620 8758 864
rect 9010 620 9016 864
rect 8752 614 9016 620
rect 9428 870 9848 876
rect 11533 870 11603 909
rect 9428 620 9440 870
rect 9836 864 10620 870
rect 9836 806 10194 864
rect 10614 806 10620 864
rect 9836 800 10620 806
rect 10770 864 11603 870
rect 10770 806 10776 864
rect 11196 806 11603 864
rect 10770 800 11603 806
rect 9836 620 9848 800
rect 9428 614 9848 620
rect 16122 463 16157 999
rect 16688 463 16722 999
rect 16122 90 16722 463
rect 11406 -326 11591 -316
rect 11406 -491 11416 -326
rect 11580 -491 11591 -326
rect 11406 -501 11591 -491
rect 11240 -1114 11646 -1104
rect 11240 -1182 11250 -1114
rect 11428 -1182 11646 -1114
rect 11240 -1192 11646 -1182
rect 13704 -2051 14611 -2007
rect 13704 -2433 13770 -2051
rect 14552 -2433 14611 -2051
rect 13704 -2478 14611 -2433
<< via2 >>
rect 4575 5954 4814 19057
rect 16726 18811 16952 19074
rect 14963 5804 15226 18450
rect 15841 16880 16441 17480
rect 17237 16880 17837 17480
rect 15453 16368 18221 16596
rect 15841 15484 16441 16084
rect 17237 15484 17837 16084
rect 15453 14972 18221 15200
rect 15841 14088 16441 14688
rect 17237 14088 17837 14688
rect 15453 13576 18221 13804
rect 15841 12692 16441 13292
rect 17237 12692 17837 13292
rect 15453 12180 18221 12408
rect 15841 11296 16441 11896
rect 17237 11296 17837 11896
rect 15453 10784 18221 11012
rect 15841 9900 16441 10500
rect 17237 9900 17837 10500
rect 15453 9388 18221 9616
rect 15841 8504 16441 9104
rect 17237 8504 17837 9104
rect 15453 7992 18221 8220
rect 15841 7108 16441 7708
rect 17237 7108 17837 7708
rect 7152 5334 12579 5493
rect 7152 5070 12579 5334
rect 5738 4878 6158 4936
rect 4508 2298 4692 2580
rect 14903 4225 15493 4815
rect 4885 4050 5003 4143
rect 4885 2166 4964 2239
rect 6452 724 7488 1345
rect 15440 1626 15836 1811
rect 10460 1164 11242 1546
rect 16157 463 16688 999
rect 11416 -491 11580 -326
rect 11250 -1182 11428 -1114
rect 13770 -2433 14552 -2051
<< metal3 >>
rect 4555 19074 16964 19086
rect 4555 19057 16726 19074
rect 4555 5954 4575 19057
rect 4814 18811 16726 19057
rect 16952 18811 16964 19074
rect 4814 18801 16964 18811
rect 4814 18322 4840 18801
rect 14832 18450 15258 18480
rect 14832 18416 14963 18450
rect 4814 18258 4920 18322
rect 4814 18006 4840 18258
rect 14929 18164 14963 18416
rect 14832 18100 14963 18164
rect 4814 17942 4920 18006
rect 4814 17690 4840 17942
rect 14929 17848 14963 18100
rect 14832 17784 14963 17848
rect 4814 17626 4920 17690
rect 4814 17374 4840 17626
rect 14929 17532 14963 17784
rect 14832 17468 14963 17532
rect 4814 17310 4920 17374
rect 4814 17058 4840 17310
rect 14929 17216 14963 17468
rect 14832 17152 14963 17216
rect 4814 16994 4920 17058
rect 4814 16742 4840 16994
rect 14929 16900 14963 17152
rect 14832 16836 14963 16900
rect 4814 16678 4920 16742
rect 4814 16426 4840 16678
rect 14929 16584 14963 16836
rect 14832 16520 14963 16584
rect 4814 16362 4920 16426
rect 4814 16110 4840 16362
rect 14929 16268 14963 16520
rect 14832 16204 14963 16268
rect 4814 16046 4920 16110
rect 4814 15794 4840 16046
rect 14929 15952 14963 16204
rect 14832 15888 14963 15952
rect 4814 15730 4920 15794
rect 4814 15478 4840 15730
rect 14929 15636 14963 15888
rect 14832 15572 14963 15636
rect 4814 15414 4920 15478
rect 4814 15162 4840 15414
rect 14929 15320 14963 15572
rect 14832 15256 14963 15320
rect 4814 15098 4920 15162
rect 4814 14846 4840 15098
rect 14929 15004 14963 15256
rect 14832 14940 14963 15004
rect 4814 14782 4920 14846
rect 4814 14530 4840 14782
rect 14929 14688 14963 14940
rect 14832 14624 14963 14688
rect 4814 14466 4920 14530
rect 4814 14214 4840 14466
rect 14929 14372 14963 14624
rect 14832 14308 14963 14372
rect 4814 14150 4920 14214
rect 4814 13898 4840 14150
rect 14929 14056 14963 14308
rect 14832 13992 14963 14056
rect 4814 13834 4920 13898
rect 4814 13582 4840 13834
rect 14929 13740 14963 13992
rect 14832 13676 14963 13740
rect 4814 13518 4920 13582
rect 4814 13266 4840 13518
rect 14929 13424 14963 13676
rect 14832 13360 14963 13424
rect 4814 13202 4920 13266
rect 4814 12950 4840 13202
rect 14929 13108 14963 13360
rect 14832 13044 14963 13108
rect 4814 12886 4920 12950
rect 4814 12634 4840 12886
rect 14929 12792 14963 13044
rect 14832 12728 14963 12792
rect 4814 12570 4920 12634
rect 4814 12318 4840 12570
rect 14929 12476 14963 12728
rect 14832 12412 14963 12476
rect 4814 12254 4920 12318
rect 4814 12002 4840 12254
rect 14929 12160 14963 12412
rect 14832 12096 14963 12160
rect 4814 11938 4920 12002
rect 4814 11686 4840 11938
rect 14929 11844 14963 12096
rect 14832 11780 14963 11844
rect 4814 11622 4920 11686
rect 4814 11370 4840 11622
rect 14929 11528 14963 11780
rect 14832 11464 14963 11528
rect 4814 11306 4920 11370
rect 4814 11054 4840 11306
rect 14929 11212 14963 11464
rect 14832 11148 14963 11212
rect 4814 10990 4920 11054
rect 4814 10738 4840 10990
rect 14929 10896 14963 11148
rect 14832 10832 14963 10896
rect 4814 10674 4920 10738
rect 4814 10422 4840 10674
rect 14929 10580 14963 10832
rect 14832 10516 14963 10580
rect 4814 10358 4920 10422
rect 4814 10106 4840 10358
rect 14929 10264 14963 10516
rect 14832 10200 14963 10264
rect 4814 10042 4920 10106
rect 4814 9790 4840 10042
rect 14929 9948 14963 10200
rect 14832 9884 14963 9948
rect 4814 9726 4920 9790
rect 4814 9474 4840 9726
rect 14929 9632 14963 9884
rect 14832 9568 14963 9632
rect 4814 9410 4920 9474
rect 4814 9158 4840 9410
rect 14929 9316 14963 9568
rect 14832 9252 14963 9316
rect 4814 9094 4920 9158
rect 4814 8842 4840 9094
rect 14929 9000 14963 9252
rect 14832 8936 14963 9000
rect 4814 8778 4920 8842
rect 4814 8526 4840 8778
rect 14929 8684 14963 8936
rect 14832 8620 14963 8684
rect 4814 8462 4920 8526
rect 4814 8210 4840 8462
rect 14929 8368 14963 8620
rect 14832 8304 14963 8368
rect 4814 8146 4920 8210
rect 4814 7894 4840 8146
rect 14929 8052 14963 8304
rect 14832 7988 14963 8052
rect 4814 7830 4920 7894
rect 4814 7578 4840 7830
rect 14929 7736 14963 7988
rect 14832 7672 14963 7736
rect 4814 7514 4920 7578
rect 4814 7262 4840 7514
rect 14929 7420 14963 7672
rect 14832 7356 14963 7420
rect 4814 7198 4920 7262
rect 4814 6946 4840 7198
rect 14929 7104 14963 7356
rect 14832 7040 14963 7104
rect 4814 6882 4920 6946
rect 4814 6630 4840 6882
rect 14929 6788 14963 7040
rect 14832 6724 14963 6788
rect 4814 6566 4920 6630
rect 4814 6314 4840 6566
rect 14929 6472 14963 6724
rect 14832 6408 14963 6472
rect 4814 6250 4920 6314
rect 4814 5998 4840 6250
rect 14929 6156 14963 6408
rect 14832 6092 14963 6156
rect 4814 5954 4920 5998
rect 4555 5934 4920 5954
rect 4555 5933 4840 5934
rect 14929 5840 14963 6092
rect 14832 5804 14963 5840
rect 15226 17480 15258 18450
rect 15741 17480 16541 17580
rect 17137 17480 17937 17580
rect 15226 16880 15841 17480
rect 16441 16880 17237 17480
rect 17837 16880 17937 17480
rect 15226 16084 15258 16880
rect 15741 16780 16541 16880
rect 17137 16780 17937 16880
rect 15443 16596 18637 16606
rect 15443 16368 15453 16596
rect 18221 16368 18637 16596
rect 15443 16358 18637 16368
rect 15741 16084 16541 16184
rect 17137 16084 17937 16184
rect 15226 15484 15841 16084
rect 16441 15484 17237 16084
rect 17837 15484 17937 16084
rect 15226 14688 15258 15484
rect 15741 15384 16541 15484
rect 17137 15384 17937 15484
rect 18463 15210 18637 16358
rect 15443 15200 18637 15210
rect 15443 14972 15453 15200
rect 18221 14972 18637 15200
rect 15443 14962 18637 14972
rect 15741 14688 16541 14788
rect 17137 14688 17937 14788
rect 15226 14088 15841 14688
rect 16441 14088 17237 14688
rect 17837 14088 17937 14688
rect 15226 13292 15258 14088
rect 15741 13988 16541 14088
rect 17137 13988 17937 14088
rect 18463 13814 18637 14962
rect 15443 13804 18637 13814
rect 15443 13576 15453 13804
rect 18221 13576 18637 13804
rect 15443 13566 18637 13576
rect 15741 13292 16541 13392
rect 17137 13292 17937 13392
rect 15226 12692 15841 13292
rect 16441 12692 17237 13292
rect 17837 12692 17937 13292
rect 15226 11896 15258 12692
rect 15741 12592 16541 12692
rect 17137 12592 17937 12692
rect 18463 12418 18637 13566
rect 15443 12408 18637 12418
rect 15443 12180 15453 12408
rect 18221 12180 18637 12408
rect 15443 12170 18637 12180
rect 15741 11896 16541 11996
rect 17137 11896 17937 11996
rect 15226 11296 15841 11896
rect 16441 11296 17237 11896
rect 17837 11296 17937 11896
rect 15226 10500 15258 11296
rect 15741 11196 16541 11296
rect 17137 11196 17937 11296
rect 18463 11022 18637 12170
rect 15443 11012 18637 11022
rect 15443 10784 15453 11012
rect 18221 10784 18637 11012
rect 15443 10774 18637 10784
rect 15741 10500 16541 10600
rect 17137 10500 17937 10600
rect 15226 9900 15841 10500
rect 16441 9900 17237 10500
rect 17837 9900 17937 10500
rect 15226 9104 15258 9900
rect 15741 9800 16541 9900
rect 17137 9800 17937 9900
rect 18463 9626 18637 10774
rect 15443 9616 18637 9626
rect 15443 9388 15453 9616
rect 18221 9388 18637 9616
rect 15443 9378 18637 9388
rect 15741 9104 16541 9204
rect 17137 9104 17937 9204
rect 15226 8504 15841 9104
rect 16441 8504 17237 9104
rect 17837 8504 17937 9104
rect 15226 7708 15258 8504
rect 15741 8404 16541 8504
rect 17137 8404 17937 8504
rect 18463 8230 18637 9378
rect 15443 8220 18637 8230
rect 15443 7992 15453 8220
rect 18221 7992 18637 8220
rect 15443 7982 18637 7992
rect 15741 7708 16541 7808
rect 17137 7708 17937 7808
rect 15226 7108 15841 7708
rect 16441 7108 17237 7708
rect 17837 7108 17937 7708
rect 15226 5804 15258 7108
rect 15741 7008 16541 7108
rect 17137 7008 17937 7108
rect 14832 5776 15258 5804
rect 7098 5493 12654 5552
rect 7098 5070 7152 5493
rect 12579 5070 12654 5493
rect 7098 5019 12654 5070
rect 5726 4936 6170 4948
rect 5726 4878 5738 4936
rect 6158 4886 6170 4936
rect 6158 4878 9644 4886
rect 5726 4774 9644 4878
rect 4876 4143 5012 4151
rect 4876 4050 4885 4143
rect 5003 4050 5012 4143
rect 9532 4091 9644 4774
rect 14898 4815 16722 4820
rect 14898 4318 14903 4815
rect 15493 4318 16722 4815
rect 4876 4043 5012 4050
rect 4498 2580 4702 2588
rect 4498 2298 4508 2580
rect 4692 2298 4702 2580
rect 4498 -56 4702 2298
rect 4876 2239 4974 4043
rect 9527 3981 9533 4091
rect 9643 3981 9649 4091
rect 9532 3980 9644 3981
rect 14894 3718 14900 4318
rect 15500 4220 16722 4318
rect 15500 3718 15506 4220
rect 4876 2166 4885 2239
rect 4964 2166 4974 2239
rect 4876 2156 4974 2166
rect 15422 1811 15854 1832
rect 15422 1626 15440 1811
rect 15836 1626 15854 1811
rect 15422 1608 15854 1626
rect 10394 1546 11301 1590
rect 6393 1345 7554 1390
rect 6393 724 6452 1345
rect 7488 724 7554 1345
rect 10394 1164 10460 1546
rect 11242 1164 11301 1546
rect 10394 1119 11301 1164
rect 6393 680 7554 724
rect 16122 999 16722 4220
rect 16122 463 16157 999
rect 16688 463 16722 999
rect 16122 434 16722 463
rect 4498 -306 4508 -56
rect 4692 -112 4702 -56
rect 4692 -306 5328 -112
rect 4498 -316 5328 -306
rect 11406 -326 11591 -316
rect 11406 -491 11416 -326
rect 11580 -491 11591 -326
rect 11406 -501 11591 -491
rect 11240 -1114 11440 -1104
rect 11240 -1182 11250 -1114
rect 11428 -1182 11440 -1114
rect 11240 -1192 11440 -1182
rect 13704 -2051 14611 -2007
rect 13704 -2433 13770 -2051
rect 14552 -2433 14611 -2051
rect 13704 -2478 14611 -2433
<< via3 >>
rect 4575 5954 4814 19057
rect 14963 5804 15226 18450
rect 7152 5070 12579 5493
rect 9533 3981 9643 4091
rect 14900 4225 14903 4318
rect 14903 4225 15493 4318
rect 15493 4225 15500 4318
rect 14900 3718 15500 4225
rect 15440 1626 15836 1811
rect 6452 724 7488 1345
rect 10460 1164 11242 1546
rect 4508 -306 4692 -56
rect 11416 -491 11580 -326
rect 11250 -1182 11428 -1114
rect 13770 -2433 14552 -2051
<< metal4 >>
rect 4555 19057 4840 19086
rect 4555 5954 4575 19057
rect 4814 5954 4840 19057
rect 4555 5933 4840 5954
rect 14929 18450 15258 18480
rect 14929 5804 14963 18450
rect 15226 5804 15258 18450
rect 14929 5776 15258 5804
rect 7098 5493 17001 5552
rect 7098 5070 7152 5493
rect 12579 5070 17001 5493
rect 7098 5019 17001 5070
rect 9532 4091 9644 4092
rect 9532 3981 9533 4091
rect 9643 3981 9644 4091
rect 9532 3518 9644 3981
rect 9532 3406 12340 3518
rect 15422 1811 15854 1832
rect 14689 1626 15440 1811
rect 15836 1626 15854 1811
rect 10394 1546 11301 1590
rect 6393 1345 7554 1390
rect 6393 724 6452 1345
rect 7488 724 7554 1345
rect 6393 680 7554 724
rect 4440 -56 4702 -46
rect 4440 -316 4454 -56
rect 4694 -316 4702 -56
rect 7908 -62 8278 1476
rect 10394 1164 10460 1546
rect 11242 1164 11301 1546
rect 10394 1119 11301 1164
rect 14689 1077 14874 1626
rect 15422 1608 15854 1626
rect 11500 892 14874 1077
rect 11500 -316 11685 892
rect 16401 178 17001 5019
rect 4440 -330 4702 -316
rect 11406 -326 11685 -316
rect 11406 -491 11416 -326
rect 11580 -491 11685 -326
rect 11406 -501 11685 -491
rect 9080 -1114 11440 -1038
rect 9080 -1182 11250 -1114
rect 11428 -1182 11440 -1114
rect 9080 -1264 11440 -1182
rect 13704 -2051 14611 -2007
rect 13704 -2433 13770 -2051
rect 14552 -2433 14611 -2051
rect 13704 -2478 14611 -2433
<< via4 >>
rect 4575 5954 4814 19057
rect 14963 5804 15226 18450
rect 14899 4318 15501 4319
rect 14899 3718 14900 4318
rect 14900 3718 15500 4318
rect 15500 3718 15501 4318
rect 14899 3717 15501 3718
rect 6452 724 7488 1345
rect 4454 -306 4508 -56
rect 4508 -306 4692 -56
rect 4692 -306 4694 -56
rect 4454 -316 4694 -306
rect 10460 1164 11242 1546
rect 13770 -2433 14552 -2051
<< metal5 >>
rect 4512 19057 4840 19086
rect 4512 5954 4575 19057
rect 4814 5954 4840 19057
rect 4512 1109 4840 5954
rect 14929 18450 15258 18703
rect 14929 5804 14963 18450
rect 15226 5804 15258 18450
rect 14929 5776 15258 5804
rect 14875 4319 15525 4343
rect 14875 3717 14899 4319
rect 15501 3717 15525 4319
rect 14875 3693 15525 3717
rect 10394 1546 11301 1590
rect 6393 1345 7554 1390
rect 6393 1109 6452 1345
rect 4512 781 6452 1109
rect 6393 724 6452 781
rect 7488 1119 7554 1345
rect 10394 1164 10460 1546
rect 11242 1164 11301 1546
rect 10394 1119 11301 1164
rect 7488 724 11301 1119
rect 6393 680 11301 724
rect 4398 -56 5134 -12
rect 4398 -316 4454 -56
rect 4694 -316 5134 -56
rect 4398 -412 5134 -316
rect 10817 -2007 11301 680
rect 10817 -2051 14611 -2007
rect 10817 -2433 13770 -2051
rect 14552 -2433 14611 -2051
rect 10817 -2478 14611 -2433
use large_nmos_g5d10  large_nmos_g5d10_0
timestamp 1664842101
transform 0 1 4986 -1 0 18582
box -124 -66 13030 4890
use large_nmos_g5d10  large_nmos_g5d10_1
timestamp 1664842101
transform 0 1 9942 -1 0 18582
box -124 -66 13030 4890
use opamp_big  opamp_big_0
timestamp 1665943203
transform 1 0 12086 0 1 -1124
box -460 -1056 5706 1930
use opamp_small  opamp_small_0
timestamp 1665942972
transform 1 0 5335 0 1 2342
box -461 -954 4014 2020
use opamp_small  opamp_small_1
timestamp 1665942972
transform 1 0 10409 0 1 2342
box -461 -954 4014 2020
use sky130_fd_pr__cap_mim_m3_1_EZNXMG  sky130_fd_pr__cap_mim_m3_1_EZNXMG_0
timestamp 1665944152
transform 1 0 7070 0 1 -1058
box -2150 -1100 2048 1100
use sky130_fd_pr__cap_mim_m3_2_EZNXMG  sky130_fd_pr__cap_mim_m3_2_EZNXMG_0
timestamp 1665944614
transform 1 0 7271 0 1 -1058
box -2351 -1100 1849 1100
use sky130_fd_pr__diode_pd2nw_11v0_N4GF4K  sky130_fd_pr__diode_pd2nw_11v0_N4GF4K_0
timestamp 1665674841
transform 1 0 16839 0 1 12294
box -1576 -5764 1576 5764
use sky130_fd_pr__res_xhigh_po_0p35_GYHWU2  sky130_fd_pr__res_xhigh_po_0p35_GYHWU2_0
timestamp 1665944838
transform 0 1 5657 -1 0 4907
box -201 -673 201 673
use sky130_fd_pr__res_xhigh_po_0p35_GYHWU2  sky130_fd_pr__res_xhigh_po_0p35_GYHWU2_1
timestamp 1665944838
transform 0 1 10695 -1 0 835
box -201 -673 201 673
use sky130_fd_pr__res_xhigh_po_0p35_X9YLXN  sky130_fd_pr__res_xhigh_po_0p35_X9YLXN_0
timestamp 1666045574
transform 0 1 15965 -1 0 1524
box -201 -709 201 709
use sky130_fd_pr__res_xhigh_po_0p35_X9YLXN  sky130_fd_pr__res_xhigh_po_0p35_X9YLXN_1
timestamp 1666045574
transform 0 1 15965 -1 0 2242
box -201 -709 201 709
use sky130_fd_pr__res_xhigh_po_1p41_YC7ZJC  sky130_fd_pr__res_xhigh_po_1p41_YC7ZJC_0
timestamp 1665944614
transform 0 1 9300 -1 0 745
box -307 -720 307 720
<< end >>
