magic
tech sky130A
magscale 1 2
timestamp 1666296061
<< nwell >>
rect -308 -82539 308 82539
<< mvpmos >>
rect -50 74242 50 82242
rect -50 66006 50 74006
rect -50 57770 50 65770
rect -50 49534 50 57534
rect -50 41298 50 49298
rect -50 33062 50 41062
rect -50 24826 50 32826
rect -50 16590 50 24590
rect -50 8354 50 16354
rect -50 118 50 8118
rect -50 -8118 50 -118
rect -50 -16354 50 -8354
rect -50 -24590 50 -16590
rect -50 -32826 50 -24826
rect -50 -41062 50 -33062
rect -50 -49298 50 -41298
rect -50 -57534 50 -49534
rect -50 -65770 50 -57770
rect -50 -74006 50 -66006
rect -50 -82242 50 -74242
<< mvpdiff >>
rect -108 82230 -50 82242
rect -108 74254 -96 82230
rect -62 74254 -50 82230
rect -108 74242 -50 74254
rect 50 82230 108 82242
rect 50 74254 62 82230
rect 96 74254 108 82230
rect 50 74242 108 74254
rect -108 73994 -50 74006
rect -108 66018 -96 73994
rect -62 66018 -50 73994
rect -108 66006 -50 66018
rect 50 73994 108 74006
rect 50 66018 62 73994
rect 96 66018 108 73994
rect 50 66006 108 66018
rect -108 65758 -50 65770
rect -108 57782 -96 65758
rect -62 57782 -50 65758
rect -108 57770 -50 57782
rect 50 65758 108 65770
rect 50 57782 62 65758
rect 96 57782 108 65758
rect 50 57770 108 57782
rect -108 57522 -50 57534
rect -108 49546 -96 57522
rect -62 49546 -50 57522
rect -108 49534 -50 49546
rect 50 57522 108 57534
rect 50 49546 62 57522
rect 96 49546 108 57522
rect 50 49534 108 49546
rect -108 49286 -50 49298
rect -108 41310 -96 49286
rect -62 41310 -50 49286
rect -108 41298 -50 41310
rect 50 49286 108 49298
rect 50 41310 62 49286
rect 96 41310 108 49286
rect 50 41298 108 41310
rect -108 41050 -50 41062
rect -108 33074 -96 41050
rect -62 33074 -50 41050
rect -108 33062 -50 33074
rect 50 41050 108 41062
rect 50 33074 62 41050
rect 96 33074 108 41050
rect 50 33062 108 33074
rect -108 32814 -50 32826
rect -108 24838 -96 32814
rect -62 24838 -50 32814
rect -108 24826 -50 24838
rect 50 32814 108 32826
rect 50 24838 62 32814
rect 96 24838 108 32814
rect 50 24826 108 24838
rect -108 24578 -50 24590
rect -108 16602 -96 24578
rect -62 16602 -50 24578
rect -108 16590 -50 16602
rect 50 24578 108 24590
rect 50 16602 62 24578
rect 96 16602 108 24578
rect 50 16590 108 16602
rect -108 16342 -50 16354
rect -108 8366 -96 16342
rect -62 8366 -50 16342
rect -108 8354 -50 8366
rect 50 16342 108 16354
rect 50 8366 62 16342
rect 96 8366 108 16342
rect 50 8354 108 8366
rect -108 8106 -50 8118
rect -108 130 -96 8106
rect -62 130 -50 8106
rect -108 118 -50 130
rect 50 8106 108 8118
rect 50 130 62 8106
rect 96 130 108 8106
rect 50 118 108 130
rect -108 -130 -50 -118
rect -108 -8106 -96 -130
rect -62 -8106 -50 -130
rect -108 -8118 -50 -8106
rect 50 -130 108 -118
rect 50 -8106 62 -130
rect 96 -8106 108 -130
rect 50 -8118 108 -8106
rect -108 -8366 -50 -8354
rect -108 -16342 -96 -8366
rect -62 -16342 -50 -8366
rect -108 -16354 -50 -16342
rect 50 -8366 108 -8354
rect 50 -16342 62 -8366
rect 96 -16342 108 -8366
rect 50 -16354 108 -16342
rect -108 -16602 -50 -16590
rect -108 -24578 -96 -16602
rect -62 -24578 -50 -16602
rect -108 -24590 -50 -24578
rect 50 -16602 108 -16590
rect 50 -24578 62 -16602
rect 96 -24578 108 -16602
rect 50 -24590 108 -24578
rect -108 -24838 -50 -24826
rect -108 -32814 -96 -24838
rect -62 -32814 -50 -24838
rect -108 -32826 -50 -32814
rect 50 -24838 108 -24826
rect 50 -32814 62 -24838
rect 96 -32814 108 -24838
rect 50 -32826 108 -32814
rect -108 -33074 -50 -33062
rect -108 -41050 -96 -33074
rect -62 -41050 -50 -33074
rect -108 -41062 -50 -41050
rect 50 -33074 108 -33062
rect 50 -41050 62 -33074
rect 96 -41050 108 -33074
rect 50 -41062 108 -41050
rect -108 -41310 -50 -41298
rect -108 -49286 -96 -41310
rect -62 -49286 -50 -41310
rect -108 -49298 -50 -49286
rect 50 -41310 108 -41298
rect 50 -49286 62 -41310
rect 96 -49286 108 -41310
rect 50 -49298 108 -49286
rect -108 -49546 -50 -49534
rect -108 -57522 -96 -49546
rect -62 -57522 -50 -49546
rect -108 -57534 -50 -57522
rect 50 -49546 108 -49534
rect 50 -57522 62 -49546
rect 96 -57522 108 -49546
rect 50 -57534 108 -57522
rect -108 -57782 -50 -57770
rect -108 -65758 -96 -57782
rect -62 -65758 -50 -57782
rect -108 -65770 -50 -65758
rect 50 -57782 108 -57770
rect 50 -65758 62 -57782
rect 96 -65758 108 -57782
rect 50 -65770 108 -65758
rect -108 -66018 -50 -66006
rect -108 -73994 -96 -66018
rect -62 -73994 -50 -66018
rect -108 -74006 -50 -73994
rect 50 -66018 108 -66006
rect 50 -73994 62 -66018
rect 96 -73994 108 -66018
rect 50 -74006 108 -73994
rect -108 -74254 -50 -74242
rect -108 -82230 -96 -74254
rect -62 -82230 -50 -74254
rect -108 -82242 -50 -82230
rect 50 -74254 108 -74242
rect 50 -82230 62 -74254
rect 96 -82230 108 -74254
rect 50 -82242 108 -82230
<< mvpdiffc >>
rect -96 74254 -62 82230
rect 62 74254 96 82230
rect -96 66018 -62 73994
rect 62 66018 96 73994
rect -96 57782 -62 65758
rect 62 57782 96 65758
rect -96 49546 -62 57522
rect 62 49546 96 57522
rect -96 41310 -62 49286
rect 62 41310 96 49286
rect -96 33074 -62 41050
rect 62 33074 96 41050
rect -96 24838 -62 32814
rect 62 24838 96 32814
rect -96 16602 -62 24578
rect 62 16602 96 24578
rect -96 8366 -62 16342
rect 62 8366 96 16342
rect -96 130 -62 8106
rect 62 130 96 8106
rect -96 -8106 -62 -130
rect 62 -8106 96 -130
rect -96 -16342 -62 -8366
rect 62 -16342 96 -8366
rect -96 -24578 -62 -16602
rect 62 -24578 96 -16602
rect -96 -32814 -62 -24838
rect 62 -32814 96 -24838
rect -96 -41050 -62 -33074
rect 62 -41050 96 -33074
rect -96 -49286 -62 -41310
rect 62 -49286 96 -41310
rect -96 -57522 -62 -49546
rect 62 -57522 96 -49546
rect -96 -65758 -62 -57782
rect 62 -65758 96 -57782
rect -96 -73994 -62 -66018
rect 62 -73994 96 -66018
rect -96 -82230 -62 -74254
rect 62 -82230 96 -74254
<< mvnsubdiff >>
rect -242 82461 242 82473
rect -242 82427 -134 82461
rect 134 82427 242 82461
rect -242 82415 242 82427
rect -242 82365 -184 82415
rect -242 -82365 -230 82365
rect -196 -82365 -184 82365
rect 184 82365 242 82415
rect -242 -82415 -184 -82365
rect 184 -82365 196 82365
rect 230 -82365 242 82365
rect 184 -82415 242 -82365
rect -242 -82427 242 -82415
rect -242 -82461 -134 -82427
rect 134 -82461 242 -82427
rect -242 -82473 242 -82461
<< mvnsubdiffcont >>
rect -134 82427 134 82461
rect -230 -82365 -196 82365
rect 196 -82365 230 82365
rect -134 -82461 134 -82427
<< poly >>
rect -50 82323 50 82339
rect -50 82289 -34 82323
rect 34 82289 50 82323
rect -50 82242 50 82289
rect -50 74195 50 74242
rect -50 74161 -34 74195
rect 34 74161 50 74195
rect -50 74145 50 74161
rect -50 74087 50 74103
rect -50 74053 -34 74087
rect 34 74053 50 74087
rect -50 74006 50 74053
rect -50 65959 50 66006
rect -50 65925 -34 65959
rect 34 65925 50 65959
rect -50 65909 50 65925
rect -50 65851 50 65867
rect -50 65817 -34 65851
rect 34 65817 50 65851
rect -50 65770 50 65817
rect -50 57723 50 57770
rect -50 57689 -34 57723
rect 34 57689 50 57723
rect -50 57673 50 57689
rect -50 57615 50 57631
rect -50 57581 -34 57615
rect 34 57581 50 57615
rect -50 57534 50 57581
rect -50 49487 50 49534
rect -50 49453 -34 49487
rect 34 49453 50 49487
rect -50 49437 50 49453
rect -50 49379 50 49395
rect -50 49345 -34 49379
rect 34 49345 50 49379
rect -50 49298 50 49345
rect -50 41251 50 41298
rect -50 41217 -34 41251
rect 34 41217 50 41251
rect -50 41201 50 41217
rect -50 41143 50 41159
rect -50 41109 -34 41143
rect 34 41109 50 41143
rect -50 41062 50 41109
rect -50 33015 50 33062
rect -50 32981 -34 33015
rect 34 32981 50 33015
rect -50 32965 50 32981
rect -50 32907 50 32923
rect -50 32873 -34 32907
rect 34 32873 50 32907
rect -50 32826 50 32873
rect -50 24779 50 24826
rect -50 24745 -34 24779
rect 34 24745 50 24779
rect -50 24729 50 24745
rect -50 24671 50 24687
rect -50 24637 -34 24671
rect 34 24637 50 24671
rect -50 24590 50 24637
rect -50 16543 50 16590
rect -50 16509 -34 16543
rect 34 16509 50 16543
rect -50 16493 50 16509
rect -50 16435 50 16451
rect -50 16401 -34 16435
rect 34 16401 50 16435
rect -50 16354 50 16401
rect -50 8307 50 8354
rect -50 8273 -34 8307
rect 34 8273 50 8307
rect -50 8257 50 8273
rect -50 8199 50 8215
rect -50 8165 -34 8199
rect 34 8165 50 8199
rect -50 8118 50 8165
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -8165 50 -8118
rect -50 -8199 -34 -8165
rect 34 -8199 50 -8165
rect -50 -8215 50 -8199
rect -50 -8273 50 -8257
rect -50 -8307 -34 -8273
rect 34 -8307 50 -8273
rect -50 -8354 50 -8307
rect -50 -16401 50 -16354
rect -50 -16435 -34 -16401
rect 34 -16435 50 -16401
rect -50 -16451 50 -16435
rect -50 -16509 50 -16493
rect -50 -16543 -34 -16509
rect 34 -16543 50 -16509
rect -50 -16590 50 -16543
rect -50 -24637 50 -24590
rect -50 -24671 -34 -24637
rect 34 -24671 50 -24637
rect -50 -24687 50 -24671
rect -50 -24745 50 -24729
rect -50 -24779 -34 -24745
rect 34 -24779 50 -24745
rect -50 -24826 50 -24779
rect -50 -32873 50 -32826
rect -50 -32907 -34 -32873
rect 34 -32907 50 -32873
rect -50 -32923 50 -32907
rect -50 -32981 50 -32965
rect -50 -33015 -34 -32981
rect 34 -33015 50 -32981
rect -50 -33062 50 -33015
rect -50 -41109 50 -41062
rect -50 -41143 -34 -41109
rect 34 -41143 50 -41109
rect -50 -41159 50 -41143
rect -50 -41217 50 -41201
rect -50 -41251 -34 -41217
rect 34 -41251 50 -41217
rect -50 -41298 50 -41251
rect -50 -49345 50 -49298
rect -50 -49379 -34 -49345
rect 34 -49379 50 -49345
rect -50 -49395 50 -49379
rect -50 -49453 50 -49437
rect -50 -49487 -34 -49453
rect 34 -49487 50 -49453
rect -50 -49534 50 -49487
rect -50 -57581 50 -57534
rect -50 -57615 -34 -57581
rect 34 -57615 50 -57581
rect -50 -57631 50 -57615
rect -50 -57689 50 -57673
rect -50 -57723 -34 -57689
rect 34 -57723 50 -57689
rect -50 -57770 50 -57723
rect -50 -65817 50 -65770
rect -50 -65851 -34 -65817
rect 34 -65851 50 -65817
rect -50 -65867 50 -65851
rect -50 -65925 50 -65909
rect -50 -65959 -34 -65925
rect 34 -65959 50 -65925
rect -50 -66006 50 -65959
rect -50 -74053 50 -74006
rect -50 -74087 -34 -74053
rect 34 -74087 50 -74053
rect -50 -74103 50 -74087
rect -50 -74161 50 -74145
rect -50 -74195 -34 -74161
rect 34 -74195 50 -74161
rect -50 -74242 50 -74195
rect -50 -82289 50 -82242
rect -50 -82323 -34 -82289
rect 34 -82323 50 -82289
rect -50 -82339 50 -82323
<< polycont >>
rect -34 82289 34 82323
rect -34 74161 34 74195
rect -34 74053 34 74087
rect -34 65925 34 65959
rect -34 65817 34 65851
rect -34 57689 34 57723
rect -34 57581 34 57615
rect -34 49453 34 49487
rect -34 49345 34 49379
rect -34 41217 34 41251
rect -34 41109 34 41143
rect -34 32981 34 33015
rect -34 32873 34 32907
rect -34 24745 34 24779
rect -34 24637 34 24671
rect -34 16509 34 16543
rect -34 16401 34 16435
rect -34 8273 34 8307
rect -34 8165 34 8199
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -8199 34 -8165
rect -34 -8307 34 -8273
rect -34 -16435 34 -16401
rect -34 -16543 34 -16509
rect -34 -24671 34 -24637
rect -34 -24779 34 -24745
rect -34 -32907 34 -32873
rect -34 -33015 34 -32981
rect -34 -41143 34 -41109
rect -34 -41251 34 -41217
rect -34 -49379 34 -49345
rect -34 -49487 34 -49453
rect -34 -57615 34 -57581
rect -34 -57723 34 -57689
rect -34 -65851 34 -65817
rect -34 -65959 34 -65925
rect -34 -74087 34 -74053
rect -34 -74195 34 -74161
rect -34 -82323 34 -82289
<< locali >>
rect -230 82427 -134 82461
rect 134 82427 230 82461
rect -230 82365 -196 82427
rect 196 82365 230 82427
rect -50 82289 -34 82323
rect 34 82289 50 82323
rect -96 82230 -62 82246
rect -96 74238 -62 74254
rect 62 82230 96 82246
rect 62 74238 96 74254
rect -50 74161 -34 74195
rect 34 74161 50 74195
rect -50 74053 -34 74087
rect 34 74053 50 74087
rect -96 73994 -62 74010
rect -96 66002 -62 66018
rect 62 73994 96 74010
rect 62 66002 96 66018
rect -50 65925 -34 65959
rect 34 65925 50 65959
rect -50 65817 -34 65851
rect 34 65817 50 65851
rect -96 65758 -62 65774
rect -96 57766 -62 57782
rect 62 65758 96 65774
rect 62 57766 96 57782
rect -50 57689 -34 57723
rect 34 57689 50 57723
rect -50 57581 -34 57615
rect 34 57581 50 57615
rect -96 57522 -62 57538
rect -96 49530 -62 49546
rect 62 57522 96 57538
rect 62 49530 96 49546
rect -50 49453 -34 49487
rect 34 49453 50 49487
rect -50 49345 -34 49379
rect 34 49345 50 49379
rect -96 49286 -62 49302
rect -96 41294 -62 41310
rect 62 49286 96 49302
rect 62 41294 96 41310
rect -50 41217 -34 41251
rect 34 41217 50 41251
rect -50 41109 -34 41143
rect 34 41109 50 41143
rect -96 41050 -62 41066
rect -96 33058 -62 33074
rect 62 41050 96 41066
rect 62 33058 96 33074
rect -50 32981 -34 33015
rect 34 32981 50 33015
rect -50 32873 -34 32907
rect 34 32873 50 32907
rect -96 32814 -62 32830
rect -96 24822 -62 24838
rect 62 32814 96 32830
rect 62 24822 96 24838
rect -50 24745 -34 24779
rect 34 24745 50 24779
rect -50 24637 -34 24671
rect 34 24637 50 24671
rect -96 24578 -62 24594
rect -96 16586 -62 16602
rect 62 24578 96 24594
rect 62 16586 96 16602
rect -50 16509 -34 16543
rect 34 16509 50 16543
rect -50 16401 -34 16435
rect 34 16401 50 16435
rect -96 16342 -62 16358
rect -96 8350 -62 8366
rect 62 16342 96 16358
rect 62 8350 96 8366
rect -50 8273 -34 8307
rect 34 8273 50 8307
rect -50 8165 -34 8199
rect 34 8165 50 8199
rect -96 8106 -62 8122
rect -96 114 -62 130
rect 62 8106 96 8122
rect 62 114 96 130
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -8122 -62 -8106
rect 62 -130 96 -114
rect 62 -8122 96 -8106
rect -50 -8199 -34 -8165
rect 34 -8199 50 -8165
rect -50 -8307 -34 -8273
rect 34 -8307 50 -8273
rect -96 -8366 -62 -8350
rect -96 -16358 -62 -16342
rect 62 -8366 96 -8350
rect 62 -16358 96 -16342
rect -50 -16435 -34 -16401
rect 34 -16435 50 -16401
rect -50 -16543 -34 -16509
rect 34 -16543 50 -16509
rect -96 -16602 -62 -16586
rect -96 -24594 -62 -24578
rect 62 -16602 96 -16586
rect 62 -24594 96 -24578
rect -50 -24671 -34 -24637
rect 34 -24671 50 -24637
rect -50 -24779 -34 -24745
rect 34 -24779 50 -24745
rect -96 -24838 -62 -24822
rect -96 -32830 -62 -32814
rect 62 -24838 96 -24822
rect 62 -32830 96 -32814
rect -50 -32907 -34 -32873
rect 34 -32907 50 -32873
rect -50 -33015 -34 -32981
rect 34 -33015 50 -32981
rect -96 -33074 -62 -33058
rect -96 -41066 -62 -41050
rect 62 -33074 96 -33058
rect 62 -41066 96 -41050
rect -50 -41143 -34 -41109
rect 34 -41143 50 -41109
rect -50 -41251 -34 -41217
rect 34 -41251 50 -41217
rect -96 -41310 -62 -41294
rect -96 -49302 -62 -49286
rect 62 -41310 96 -41294
rect 62 -49302 96 -49286
rect -50 -49379 -34 -49345
rect 34 -49379 50 -49345
rect -50 -49487 -34 -49453
rect 34 -49487 50 -49453
rect -96 -49546 -62 -49530
rect -96 -57538 -62 -57522
rect 62 -49546 96 -49530
rect 62 -57538 96 -57522
rect -50 -57615 -34 -57581
rect 34 -57615 50 -57581
rect -50 -57723 -34 -57689
rect 34 -57723 50 -57689
rect -96 -57782 -62 -57766
rect -96 -65774 -62 -65758
rect 62 -57782 96 -57766
rect 62 -65774 96 -65758
rect -50 -65851 -34 -65817
rect 34 -65851 50 -65817
rect -50 -65959 -34 -65925
rect 34 -65959 50 -65925
rect -96 -66018 -62 -66002
rect -96 -74010 -62 -73994
rect 62 -66018 96 -66002
rect 62 -74010 96 -73994
rect -50 -74087 -34 -74053
rect 34 -74087 50 -74053
rect -50 -74195 -34 -74161
rect 34 -74195 50 -74161
rect -96 -74254 -62 -74238
rect -96 -82246 -62 -82230
rect 62 -74254 96 -74238
rect 62 -82246 96 -82230
rect -50 -82323 -34 -82289
rect 34 -82323 50 -82289
rect -230 -82427 -196 -82365
rect 196 -82427 230 -82365
rect -230 -82461 -134 -82427
rect 134 -82461 230 -82427
<< viali >>
rect -34 82289 34 82323
rect -96 74254 -62 82230
rect 62 74254 96 82230
rect -34 74161 34 74195
rect -34 74053 34 74087
rect -96 66018 -62 73994
rect 62 66018 96 73994
rect -34 65925 34 65959
rect -34 65817 34 65851
rect -96 57782 -62 65758
rect 62 57782 96 65758
rect -34 57689 34 57723
rect -34 57581 34 57615
rect -96 49546 -62 57522
rect 62 49546 96 57522
rect -34 49453 34 49487
rect -34 49345 34 49379
rect -96 41310 -62 49286
rect 62 41310 96 49286
rect -34 41217 34 41251
rect -34 41109 34 41143
rect -96 33074 -62 41050
rect 62 33074 96 41050
rect -34 32981 34 33015
rect -34 32873 34 32907
rect -96 24838 -62 32814
rect 62 24838 96 32814
rect -34 24745 34 24779
rect -34 24637 34 24671
rect -96 16602 -62 24578
rect 62 16602 96 24578
rect -34 16509 34 16543
rect -34 16401 34 16435
rect -96 8366 -62 16342
rect 62 8366 96 16342
rect -34 8273 34 8307
rect -34 8165 34 8199
rect -96 130 -62 8106
rect 62 130 96 8106
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -8106 -62 -130
rect 62 -8106 96 -130
rect -34 -8199 34 -8165
rect -34 -8307 34 -8273
rect -96 -16342 -62 -8366
rect 62 -16342 96 -8366
rect -34 -16435 34 -16401
rect -34 -16543 34 -16509
rect -96 -24578 -62 -16602
rect 62 -24578 96 -16602
rect -34 -24671 34 -24637
rect -34 -24779 34 -24745
rect -96 -32814 -62 -24838
rect 62 -32814 96 -24838
rect -34 -32907 34 -32873
rect -34 -33015 34 -32981
rect -96 -41050 -62 -33074
rect 62 -41050 96 -33074
rect -34 -41143 34 -41109
rect -34 -41251 34 -41217
rect -96 -49286 -62 -41310
rect 62 -49286 96 -41310
rect -34 -49379 34 -49345
rect -34 -49487 34 -49453
rect -96 -57522 -62 -49546
rect 62 -57522 96 -49546
rect -34 -57615 34 -57581
rect -34 -57723 34 -57689
rect -96 -65758 -62 -57782
rect 62 -65758 96 -57782
rect -34 -65851 34 -65817
rect -34 -65959 34 -65925
rect -96 -73994 -62 -66018
rect 62 -73994 96 -66018
rect -34 -74087 34 -74053
rect -34 -74195 34 -74161
rect -96 -82230 -62 -74254
rect 62 -82230 96 -74254
rect -34 -82323 34 -82289
<< metal1 >>
rect -46 82323 46 82329
rect -46 82289 -34 82323
rect 34 82289 46 82323
rect -46 82283 46 82289
rect -102 82230 -56 82242
rect -102 74254 -96 82230
rect -62 74254 -56 82230
rect -102 74242 -56 74254
rect 56 82230 102 82242
rect 56 74254 62 82230
rect 96 74254 102 82230
rect 56 74242 102 74254
rect -46 74195 46 74201
rect -46 74161 -34 74195
rect 34 74161 46 74195
rect -46 74155 46 74161
rect -46 74087 46 74093
rect -46 74053 -34 74087
rect 34 74053 46 74087
rect -46 74047 46 74053
rect -102 73994 -56 74006
rect -102 66018 -96 73994
rect -62 66018 -56 73994
rect -102 66006 -56 66018
rect 56 73994 102 74006
rect 56 66018 62 73994
rect 96 66018 102 73994
rect 56 66006 102 66018
rect -46 65959 46 65965
rect -46 65925 -34 65959
rect 34 65925 46 65959
rect -46 65919 46 65925
rect -46 65851 46 65857
rect -46 65817 -34 65851
rect 34 65817 46 65851
rect -46 65811 46 65817
rect -102 65758 -56 65770
rect -102 57782 -96 65758
rect -62 57782 -56 65758
rect -102 57770 -56 57782
rect 56 65758 102 65770
rect 56 57782 62 65758
rect 96 57782 102 65758
rect 56 57770 102 57782
rect -46 57723 46 57729
rect -46 57689 -34 57723
rect 34 57689 46 57723
rect -46 57683 46 57689
rect -46 57615 46 57621
rect -46 57581 -34 57615
rect 34 57581 46 57615
rect -46 57575 46 57581
rect -102 57522 -56 57534
rect -102 49546 -96 57522
rect -62 49546 -56 57522
rect -102 49534 -56 49546
rect 56 57522 102 57534
rect 56 49546 62 57522
rect 96 49546 102 57522
rect 56 49534 102 49546
rect -46 49487 46 49493
rect -46 49453 -34 49487
rect 34 49453 46 49487
rect -46 49447 46 49453
rect -46 49379 46 49385
rect -46 49345 -34 49379
rect 34 49345 46 49379
rect -46 49339 46 49345
rect -102 49286 -56 49298
rect -102 41310 -96 49286
rect -62 41310 -56 49286
rect -102 41298 -56 41310
rect 56 49286 102 49298
rect 56 41310 62 49286
rect 96 41310 102 49286
rect 56 41298 102 41310
rect -46 41251 46 41257
rect -46 41217 -34 41251
rect 34 41217 46 41251
rect -46 41211 46 41217
rect -46 41143 46 41149
rect -46 41109 -34 41143
rect 34 41109 46 41143
rect -46 41103 46 41109
rect -102 41050 -56 41062
rect -102 33074 -96 41050
rect -62 33074 -56 41050
rect -102 33062 -56 33074
rect 56 41050 102 41062
rect 56 33074 62 41050
rect 96 33074 102 41050
rect 56 33062 102 33074
rect -46 33015 46 33021
rect -46 32981 -34 33015
rect 34 32981 46 33015
rect -46 32975 46 32981
rect -46 32907 46 32913
rect -46 32873 -34 32907
rect 34 32873 46 32907
rect -46 32867 46 32873
rect -102 32814 -56 32826
rect -102 24838 -96 32814
rect -62 24838 -56 32814
rect -102 24826 -56 24838
rect 56 32814 102 32826
rect 56 24838 62 32814
rect 96 24838 102 32814
rect 56 24826 102 24838
rect -46 24779 46 24785
rect -46 24745 -34 24779
rect 34 24745 46 24779
rect -46 24739 46 24745
rect -46 24671 46 24677
rect -46 24637 -34 24671
rect 34 24637 46 24671
rect -46 24631 46 24637
rect -102 24578 -56 24590
rect -102 16602 -96 24578
rect -62 16602 -56 24578
rect -102 16590 -56 16602
rect 56 24578 102 24590
rect 56 16602 62 24578
rect 96 16602 102 24578
rect 56 16590 102 16602
rect -46 16543 46 16549
rect -46 16509 -34 16543
rect 34 16509 46 16543
rect -46 16503 46 16509
rect -46 16435 46 16441
rect -46 16401 -34 16435
rect 34 16401 46 16435
rect -46 16395 46 16401
rect -102 16342 -56 16354
rect -102 8366 -96 16342
rect -62 8366 -56 16342
rect -102 8354 -56 8366
rect 56 16342 102 16354
rect 56 8366 62 16342
rect 96 8366 102 16342
rect 56 8354 102 8366
rect -46 8307 46 8313
rect -46 8273 -34 8307
rect 34 8273 46 8307
rect -46 8267 46 8273
rect -46 8199 46 8205
rect -46 8165 -34 8199
rect 34 8165 46 8199
rect -46 8159 46 8165
rect -102 8106 -56 8118
rect -102 130 -96 8106
rect -62 130 -56 8106
rect -102 118 -56 130
rect 56 8106 102 8118
rect 56 130 62 8106
rect 96 130 102 8106
rect 56 118 102 130
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -130 -56 -118
rect -102 -8106 -96 -130
rect -62 -8106 -56 -130
rect -102 -8118 -56 -8106
rect 56 -130 102 -118
rect 56 -8106 62 -130
rect 96 -8106 102 -130
rect 56 -8118 102 -8106
rect -46 -8165 46 -8159
rect -46 -8199 -34 -8165
rect 34 -8199 46 -8165
rect -46 -8205 46 -8199
rect -46 -8273 46 -8267
rect -46 -8307 -34 -8273
rect 34 -8307 46 -8273
rect -46 -8313 46 -8307
rect -102 -8366 -56 -8354
rect -102 -16342 -96 -8366
rect -62 -16342 -56 -8366
rect -102 -16354 -56 -16342
rect 56 -8366 102 -8354
rect 56 -16342 62 -8366
rect 96 -16342 102 -8366
rect 56 -16354 102 -16342
rect -46 -16401 46 -16395
rect -46 -16435 -34 -16401
rect 34 -16435 46 -16401
rect -46 -16441 46 -16435
rect -46 -16509 46 -16503
rect -46 -16543 -34 -16509
rect 34 -16543 46 -16509
rect -46 -16549 46 -16543
rect -102 -16602 -56 -16590
rect -102 -24578 -96 -16602
rect -62 -24578 -56 -16602
rect -102 -24590 -56 -24578
rect 56 -16602 102 -16590
rect 56 -24578 62 -16602
rect 96 -24578 102 -16602
rect 56 -24590 102 -24578
rect -46 -24637 46 -24631
rect -46 -24671 -34 -24637
rect 34 -24671 46 -24637
rect -46 -24677 46 -24671
rect -46 -24745 46 -24739
rect -46 -24779 -34 -24745
rect 34 -24779 46 -24745
rect -46 -24785 46 -24779
rect -102 -24838 -56 -24826
rect -102 -32814 -96 -24838
rect -62 -32814 -56 -24838
rect -102 -32826 -56 -32814
rect 56 -24838 102 -24826
rect 56 -32814 62 -24838
rect 96 -32814 102 -24838
rect 56 -32826 102 -32814
rect -46 -32873 46 -32867
rect -46 -32907 -34 -32873
rect 34 -32907 46 -32873
rect -46 -32913 46 -32907
rect -46 -32981 46 -32975
rect -46 -33015 -34 -32981
rect 34 -33015 46 -32981
rect -46 -33021 46 -33015
rect -102 -33074 -56 -33062
rect -102 -41050 -96 -33074
rect -62 -41050 -56 -33074
rect -102 -41062 -56 -41050
rect 56 -33074 102 -33062
rect 56 -41050 62 -33074
rect 96 -41050 102 -33074
rect 56 -41062 102 -41050
rect -46 -41109 46 -41103
rect -46 -41143 -34 -41109
rect 34 -41143 46 -41109
rect -46 -41149 46 -41143
rect -46 -41217 46 -41211
rect -46 -41251 -34 -41217
rect 34 -41251 46 -41217
rect -46 -41257 46 -41251
rect -102 -41310 -56 -41298
rect -102 -49286 -96 -41310
rect -62 -49286 -56 -41310
rect -102 -49298 -56 -49286
rect 56 -41310 102 -41298
rect 56 -49286 62 -41310
rect 96 -49286 102 -41310
rect 56 -49298 102 -49286
rect -46 -49345 46 -49339
rect -46 -49379 -34 -49345
rect 34 -49379 46 -49345
rect -46 -49385 46 -49379
rect -46 -49453 46 -49447
rect -46 -49487 -34 -49453
rect 34 -49487 46 -49453
rect -46 -49493 46 -49487
rect -102 -49546 -56 -49534
rect -102 -57522 -96 -49546
rect -62 -57522 -56 -49546
rect -102 -57534 -56 -57522
rect 56 -49546 102 -49534
rect 56 -57522 62 -49546
rect 96 -57522 102 -49546
rect 56 -57534 102 -57522
rect -46 -57581 46 -57575
rect -46 -57615 -34 -57581
rect 34 -57615 46 -57581
rect -46 -57621 46 -57615
rect -46 -57689 46 -57683
rect -46 -57723 -34 -57689
rect 34 -57723 46 -57689
rect -46 -57729 46 -57723
rect -102 -57782 -56 -57770
rect -102 -65758 -96 -57782
rect -62 -65758 -56 -57782
rect -102 -65770 -56 -65758
rect 56 -57782 102 -57770
rect 56 -65758 62 -57782
rect 96 -65758 102 -57782
rect 56 -65770 102 -65758
rect -46 -65817 46 -65811
rect -46 -65851 -34 -65817
rect 34 -65851 46 -65817
rect -46 -65857 46 -65851
rect -46 -65925 46 -65919
rect -46 -65959 -34 -65925
rect 34 -65959 46 -65925
rect -46 -65965 46 -65959
rect -102 -66018 -56 -66006
rect -102 -73994 -96 -66018
rect -62 -73994 -56 -66018
rect -102 -74006 -56 -73994
rect 56 -66018 102 -66006
rect 56 -73994 62 -66018
rect 96 -73994 102 -66018
rect 56 -74006 102 -73994
rect -46 -74053 46 -74047
rect -46 -74087 -34 -74053
rect 34 -74087 46 -74053
rect -46 -74093 46 -74087
rect -46 -74161 46 -74155
rect -46 -74195 -34 -74161
rect 34 -74195 46 -74161
rect -46 -74201 46 -74195
rect -102 -74254 -56 -74242
rect -102 -82230 -96 -74254
rect -62 -82230 -56 -74254
rect -102 -82242 -56 -82230
rect 56 -74254 102 -74242
rect 56 -82230 62 -74254
rect 96 -82230 102 -74254
rect 56 -82242 102 -82230
rect -46 -82289 46 -82283
rect -46 -82323 -34 -82289
rect 34 -82323 46 -82289
rect -46 -82329 46 -82323
<< properties >>
string FIXED_BBOX -213 -82444 213 82444
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 40 l 0.5 m 20 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
