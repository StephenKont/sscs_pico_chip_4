magic
tech sky130A
magscale 1 2
timestamp 1667066906
<< metal3 >>
rect -102 100750 2 100800
rect -3150 97702 3050 100750
rect -3200 97598 3100 97702
rect -3150 94550 3050 97598
rect -102 94450 2 94550
rect -3150 91402 3050 94450
rect -3200 91298 3100 91402
rect -3150 88250 3050 91298
rect -102 88150 2 88250
rect -3150 85102 3050 88150
rect -3200 84998 3100 85102
rect -3150 81950 3050 84998
rect -102 81850 2 81950
rect -3150 78802 3050 81850
rect -3200 78698 3100 78802
rect -3150 75650 3050 78698
rect -102 75550 2 75650
rect -3150 72502 3050 75550
rect -3200 72398 3100 72502
rect -3150 69350 3050 72398
rect -102 69250 2 69350
rect -3150 66202 3050 69250
rect -3200 66098 3100 66202
rect -3150 63050 3050 66098
rect -102 62950 2 63050
rect -3150 59902 3050 62950
rect -3200 59798 3100 59902
rect -3150 56750 3050 59798
rect -102 56650 2 56750
rect -3150 53602 3050 56650
rect -3200 53498 3100 53602
rect -3150 50450 3050 53498
rect -102 50350 2 50450
rect -3150 47302 3050 50350
rect -3200 47198 3100 47302
rect -3150 44150 3050 47198
rect -102 44050 2 44150
rect -3150 41002 3050 44050
rect -3200 40898 3100 41002
rect -3150 37850 3050 40898
rect -102 37750 2 37850
rect -3150 34702 3050 37750
rect -3200 34598 3100 34702
rect -3150 31550 3050 34598
rect -102 31450 2 31550
rect -3150 28402 3050 31450
rect -3200 28298 3100 28402
rect -3150 25250 3050 28298
rect -102 25150 2 25250
rect -3150 22102 3050 25150
rect -3200 21998 3100 22102
rect -3150 18950 3050 21998
rect -102 18850 2 18950
rect -3150 15802 3050 18850
rect -3200 15698 3100 15802
rect -3150 12650 3050 15698
rect -102 12550 2 12650
rect -3150 9502 3050 12550
rect -3200 9398 3100 9502
rect -3150 6350 3050 9398
rect -102 6250 2 6350
rect -3150 3202 3050 6250
rect -3200 3098 3100 3202
rect -3150 50 3050 3098
rect -102 -50 2 50
rect -3150 -3098 3050 -50
rect -3200 -3202 3100 -3098
rect -3150 -6250 3050 -3202
rect -102 -6350 2 -6250
rect -3150 -9398 3050 -6350
rect -3200 -9502 3100 -9398
rect -3150 -12550 3050 -9502
rect -102 -12650 2 -12550
rect -3150 -15698 3050 -12650
rect -3200 -15802 3100 -15698
rect -3150 -18850 3050 -15802
rect -102 -18950 2 -18850
rect -3150 -21998 3050 -18950
rect -3200 -22102 3100 -21998
rect -3150 -25150 3050 -22102
rect -102 -25250 2 -25150
rect -3150 -28298 3050 -25250
rect -3200 -28402 3100 -28298
rect -3150 -31450 3050 -28402
rect -102 -31550 2 -31450
rect -3150 -34598 3050 -31550
rect -3200 -34702 3100 -34598
rect -3150 -37750 3050 -34702
rect -102 -37850 2 -37750
rect -3150 -40898 3050 -37850
rect -3200 -41002 3100 -40898
rect -3150 -44050 3050 -41002
rect -102 -44150 2 -44050
rect -3150 -47198 3050 -44150
rect -3200 -47302 3100 -47198
rect -3150 -50350 3050 -47302
rect -102 -50450 2 -50350
rect -3150 -53498 3050 -50450
rect -3200 -53602 3100 -53498
rect -3150 -56650 3050 -53602
rect -102 -56750 2 -56650
rect -3150 -59798 3050 -56750
rect -3200 -59902 3100 -59798
rect -3150 -62950 3050 -59902
rect -102 -63050 2 -62950
rect -3150 -66098 3050 -63050
rect -3200 -66202 3100 -66098
rect -3150 -69250 3050 -66202
rect -102 -69350 2 -69250
rect -3150 -72398 3050 -69350
rect -3200 -72502 3100 -72398
rect -3150 -75550 3050 -72502
rect -102 -75650 2 -75550
rect -3150 -78698 3050 -75650
rect -3200 -78802 3100 -78698
rect -3150 -81850 3050 -78802
rect -102 -81950 2 -81850
rect -3150 -84998 3050 -81950
rect -3200 -85102 3100 -84998
rect -3150 -88150 3050 -85102
rect -102 -88250 2 -88150
rect -3150 -91298 3050 -88250
rect -3200 -91402 3100 -91298
rect -3150 -94450 3050 -91402
rect -102 -94550 2 -94450
rect -3150 -97598 3050 -94550
rect -3200 -97702 3100 -97598
rect -3150 -100750 3050 -97702
rect -102 -100800 2 -100750
<< mimcap >>
rect -3050 100610 2950 100650
rect -3050 94690 -3010 100610
rect 2910 94690 2950 100610
rect -3050 94650 2950 94690
rect -3050 94310 2950 94350
rect -3050 88390 -3010 94310
rect 2910 88390 2950 94310
rect -3050 88350 2950 88390
rect -3050 88010 2950 88050
rect -3050 82090 -3010 88010
rect 2910 82090 2950 88010
rect -3050 82050 2950 82090
rect -3050 81710 2950 81750
rect -3050 75790 -3010 81710
rect 2910 75790 2950 81710
rect -3050 75750 2950 75790
rect -3050 75410 2950 75450
rect -3050 69490 -3010 75410
rect 2910 69490 2950 75410
rect -3050 69450 2950 69490
rect -3050 69110 2950 69150
rect -3050 63190 -3010 69110
rect 2910 63190 2950 69110
rect -3050 63150 2950 63190
rect -3050 62810 2950 62850
rect -3050 56890 -3010 62810
rect 2910 56890 2950 62810
rect -3050 56850 2950 56890
rect -3050 56510 2950 56550
rect -3050 50590 -3010 56510
rect 2910 50590 2950 56510
rect -3050 50550 2950 50590
rect -3050 50210 2950 50250
rect -3050 44290 -3010 50210
rect 2910 44290 2950 50210
rect -3050 44250 2950 44290
rect -3050 43910 2950 43950
rect -3050 37990 -3010 43910
rect 2910 37990 2950 43910
rect -3050 37950 2950 37990
rect -3050 37610 2950 37650
rect -3050 31690 -3010 37610
rect 2910 31690 2950 37610
rect -3050 31650 2950 31690
rect -3050 31310 2950 31350
rect -3050 25390 -3010 31310
rect 2910 25390 2950 31310
rect -3050 25350 2950 25390
rect -3050 25010 2950 25050
rect -3050 19090 -3010 25010
rect 2910 19090 2950 25010
rect -3050 19050 2950 19090
rect -3050 18710 2950 18750
rect -3050 12790 -3010 18710
rect 2910 12790 2950 18710
rect -3050 12750 2950 12790
rect -3050 12410 2950 12450
rect -3050 6490 -3010 12410
rect 2910 6490 2950 12410
rect -3050 6450 2950 6490
rect -3050 6110 2950 6150
rect -3050 190 -3010 6110
rect 2910 190 2950 6110
rect -3050 150 2950 190
rect -3050 -190 2950 -150
rect -3050 -6110 -3010 -190
rect 2910 -6110 2950 -190
rect -3050 -6150 2950 -6110
rect -3050 -6490 2950 -6450
rect -3050 -12410 -3010 -6490
rect 2910 -12410 2950 -6490
rect -3050 -12450 2950 -12410
rect -3050 -12790 2950 -12750
rect -3050 -18710 -3010 -12790
rect 2910 -18710 2950 -12790
rect -3050 -18750 2950 -18710
rect -3050 -19090 2950 -19050
rect -3050 -25010 -3010 -19090
rect 2910 -25010 2950 -19090
rect -3050 -25050 2950 -25010
rect -3050 -25390 2950 -25350
rect -3050 -31310 -3010 -25390
rect 2910 -31310 2950 -25390
rect -3050 -31350 2950 -31310
rect -3050 -31690 2950 -31650
rect -3050 -37610 -3010 -31690
rect 2910 -37610 2950 -31690
rect -3050 -37650 2950 -37610
rect -3050 -37990 2950 -37950
rect -3050 -43910 -3010 -37990
rect 2910 -43910 2950 -37990
rect -3050 -43950 2950 -43910
rect -3050 -44290 2950 -44250
rect -3050 -50210 -3010 -44290
rect 2910 -50210 2950 -44290
rect -3050 -50250 2950 -50210
rect -3050 -50590 2950 -50550
rect -3050 -56510 -3010 -50590
rect 2910 -56510 2950 -50590
rect -3050 -56550 2950 -56510
rect -3050 -56890 2950 -56850
rect -3050 -62810 -3010 -56890
rect 2910 -62810 2950 -56890
rect -3050 -62850 2950 -62810
rect -3050 -63190 2950 -63150
rect -3050 -69110 -3010 -63190
rect 2910 -69110 2950 -63190
rect -3050 -69150 2950 -69110
rect -3050 -69490 2950 -69450
rect -3050 -75410 -3010 -69490
rect 2910 -75410 2950 -69490
rect -3050 -75450 2950 -75410
rect -3050 -75790 2950 -75750
rect -3050 -81710 -3010 -75790
rect 2910 -81710 2950 -75790
rect -3050 -81750 2950 -81710
rect -3050 -82090 2950 -82050
rect -3050 -88010 -3010 -82090
rect 2910 -88010 2950 -82090
rect -3050 -88050 2950 -88010
rect -3050 -88390 2950 -88350
rect -3050 -94310 -3010 -88390
rect 2910 -94310 2950 -88390
rect -3050 -94350 2950 -94310
rect -3050 -94690 2950 -94650
rect -3050 -100610 -3010 -94690
rect 2910 -100610 2950 -94690
rect -3050 -100650 2950 -100610
<< mimcapcontact >>
rect -3010 94690 2910 100610
rect -3010 88390 2910 94310
rect -3010 82090 2910 88010
rect -3010 75790 2910 81710
rect -3010 69490 2910 75410
rect -3010 63190 2910 69110
rect -3010 56890 2910 62810
rect -3010 50590 2910 56510
rect -3010 44290 2910 50210
rect -3010 37990 2910 43910
rect -3010 31690 2910 37610
rect -3010 25390 2910 31310
rect -3010 19090 2910 25010
rect -3010 12790 2910 18710
rect -3010 6490 2910 12410
rect -3010 190 2910 6110
rect -3010 -6110 2910 -190
rect -3010 -12410 2910 -6490
rect -3010 -18710 2910 -12790
rect -3010 -25010 2910 -19090
rect -3010 -31310 2910 -25390
rect -3010 -37610 2910 -31690
rect -3010 -43910 2910 -37990
rect -3010 -50210 2910 -44290
rect -3010 -56510 2910 -50590
rect -3010 -62810 2910 -56890
rect -3010 -69110 2910 -63190
rect -3010 -75410 2910 -69490
rect -3010 -81710 2910 -75790
rect -3010 -88010 2910 -82090
rect -3010 -94310 2910 -88390
rect -3010 -100610 2910 -94690
<< metal4 >>
rect -102 100611 2 100800
rect -3011 100610 2911 100611
rect -3011 97702 -3010 100610
rect -3200 97598 -3010 97702
rect -3011 94690 -3010 97598
rect 2910 97702 2911 100610
rect 2910 97598 3100 97702
rect 2910 94690 2911 97598
rect -3011 94689 2911 94690
rect -102 94311 2 94689
rect -3011 94310 2911 94311
rect -3011 91402 -3010 94310
rect -3200 91298 -3010 91402
rect -3011 88390 -3010 91298
rect 2910 91402 2911 94310
rect 2910 91298 3100 91402
rect 2910 88390 2911 91298
rect -3011 88389 2911 88390
rect -102 88011 2 88389
rect -3011 88010 2911 88011
rect -3011 85102 -3010 88010
rect -3200 84998 -3010 85102
rect -3011 82090 -3010 84998
rect 2910 85102 2911 88010
rect 2910 84998 3100 85102
rect 2910 82090 2911 84998
rect -3011 82089 2911 82090
rect -102 81711 2 82089
rect -3011 81710 2911 81711
rect -3011 78802 -3010 81710
rect -3200 78698 -3010 78802
rect -3011 75790 -3010 78698
rect 2910 78802 2911 81710
rect 2910 78698 3100 78802
rect 2910 75790 2911 78698
rect -3011 75789 2911 75790
rect -102 75411 2 75789
rect -3011 75410 2911 75411
rect -3011 72502 -3010 75410
rect -3200 72398 -3010 72502
rect -3011 69490 -3010 72398
rect 2910 72502 2911 75410
rect 2910 72398 3100 72502
rect 2910 69490 2911 72398
rect -3011 69489 2911 69490
rect -102 69111 2 69489
rect -3011 69110 2911 69111
rect -3011 66202 -3010 69110
rect -3200 66098 -3010 66202
rect -3011 63190 -3010 66098
rect 2910 66202 2911 69110
rect 2910 66098 3100 66202
rect 2910 63190 2911 66098
rect -3011 63189 2911 63190
rect -102 62811 2 63189
rect -3011 62810 2911 62811
rect -3011 59902 -3010 62810
rect -3200 59798 -3010 59902
rect -3011 56890 -3010 59798
rect 2910 59902 2911 62810
rect 2910 59798 3100 59902
rect 2910 56890 2911 59798
rect -3011 56889 2911 56890
rect -102 56511 2 56889
rect -3011 56510 2911 56511
rect -3011 53602 -3010 56510
rect -3200 53498 -3010 53602
rect -3011 50590 -3010 53498
rect 2910 53602 2911 56510
rect 2910 53498 3100 53602
rect 2910 50590 2911 53498
rect -3011 50589 2911 50590
rect -102 50211 2 50589
rect -3011 50210 2911 50211
rect -3011 47302 -3010 50210
rect -3200 47198 -3010 47302
rect -3011 44290 -3010 47198
rect 2910 47302 2911 50210
rect 2910 47198 3100 47302
rect 2910 44290 2911 47198
rect -3011 44289 2911 44290
rect -102 43911 2 44289
rect -3011 43910 2911 43911
rect -3011 41002 -3010 43910
rect -3200 40898 -3010 41002
rect -3011 37990 -3010 40898
rect 2910 41002 2911 43910
rect 2910 40898 3100 41002
rect 2910 37990 2911 40898
rect -3011 37989 2911 37990
rect -102 37611 2 37989
rect -3011 37610 2911 37611
rect -3011 34702 -3010 37610
rect -3200 34598 -3010 34702
rect -3011 31690 -3010 34598
rect 2910 34702 2911 37610
rect 2910 34598 3100 34702
rect 2910 31690 2911 34598
rect -3011 31689 2911 31690
rect -102 31311 2 31689
rect -3011 31310 2911 31311
rect -3011 28402 -3010 31310
rect -3200 28298 -3010 28402
rect -3011 25390 -3010 28298
rect 2910 28402 2911 31310
rect 2910 28298 3100 28402
rect 2910 25390 2911 28298
rect -3011 25389 2911 25390
rect -102 25011 2 25389
rect -3011 25010 2911 25011
rect -3011 22102 -3010 25010
rect -3200 21998 -3010 22102
rect -3011 19090 -3010 21998
rect 2910 22102 2911 25010
rect 2910 21998 3100 22102
rect 2910 19090 2911 21998
rect -3011 19089 2911 19090
rect -102 18711 2 19089
rect -3011 18710 2911 18711
rect -3011 15802 -3010 18710
rect -3200 15698 -3010 15802
rect -3011 12790 -3010 15698
rect 2910 15802 2911 18710
rect 2910 15698 3100 15802
rect 2910 12790 2911 15698
rect -3011 12789 2911 12790
rect -102 12411 2 12789
rect -3011 12410 2911 12411
rect -3011 9502 -3010 12410
rect -3200 9398 -3010 9502
rect -3011 6490 -3010 9398
rect 2910 9502 2911 12410
rect 2910 9398 3100 9502
rect 2910 6490 2911 9398
rect -3011 6489 2911 6490
rect -102 6111 2 6489
rect -3011 6110 2911 6111
rect -3011 3202 -3010 6110
rect -3200 3098 -3010 3202
rect -3011 190 -3010 3098
rect 2910 3202 2911 6110
rect 2910 3098 3100 3202
rect 2910 190 2911 3098
rect -3011 189 2911 190
rect -102 -189 2 189
rect -3011 -190 2911 -189
rect -3011 -3098 -3010 -190
rect -3200 -3202 -3010 -3098
rect -3011 -6110 -3010 -3202
rect 2910 -3098 2911 -190
rect 2910 -3202 3100 -3098
rect 2910 -6110 2911 -3202
rect -3011 -6111 2911 -6110
rect -102 -6489 2 -6111
rect -3011 -6490 2911 -6489
rect -3011 -9398 -3010 -6490
rect -3200 -9502 -3010 -9398
rect -3011 -12410 -3010 -9502
rect 2910 -9398 2911 -6490
rect 2910 -9502 3100 -9398
rect 2910 -12410 2911 -9502
rect -3011 -12411 2911 -12410
rect -102 -12789 2 -12411
rect -3011 -12790 2911 -12789
rect -3011 -15698 -3010 -12790
rect -3200 -15802 -3010 -15698
rect -3011 -18710 -3010 -15802
rect 2910 -15698 2911 -12790
rect 2910 -15802 3100 -15698
rect 2910 -18710 2911 -15802
rect -3011 -18711 2911 -18710
rect -102 -19089 2 -18711
rect -3011 -19090 2911 -19089
rect -3011 -21998 -3010 -19090
rect -3200 -22102 -3010 -21998
rect -3011 -25010 -3010 -22102
rect 2910 -21998 2911 -19090
rect 2910 -22102 3100 -21998
rect 2910 -25010 2911 -22102
rect -3011 -25011 2911 -25010
rect -102 -25389 2 -25011
rect -3011 -25390 2911 -25389
rect -3011 -28298 -3010 -25390
rect -3200 -28402 -3010 -28298
rect -3011 -31310 -3010 -28402
rect 2910 -28298 2911 -25390
rect 2910 -28402 3100 -28298
rect 2910 -31310 2911 -28402
rect -3011 -31311 2911 -31310
rect -102 -31689 2 -31311
rect -3011 -31690 2911 -31689
rect -3011 -34598 -3010 -31690
rect -3200 -34702 -3010 -34598
rect -3011 -37610 -3010 -34702
rect 2910 -34598 2911 -31690
rect 2910 -34702 3100 -34598
rect 2910 -37610 2911 -34702
rect -3011 -37611 2911 -37610
rect -102 -37989 2 -37611
rect -3011 -37990 2911 -37989
rect -3011 -40898 -3010 -37990
rect -3200 -41002 -3010 -40898
rect -3011 -43910 -3010 -41002
rect 2910 -40898 2911 -37990
rect 2910 -41002 3100 -40898
rect 2910 -43910 2911 -41002
rect -3011 -43911 2911 -43910
rect -102 -44289 2 -43911
rect -3011 -44290 2911 -44289
rect -3011 -47198 -3010 -44290
rect -3200 -47302 -3010 -47198
rect -3011 -50210 -3010 -47302
rect 2910 -47198 2911 -44290
rect 2910 -47302 3100 -47198
rect 2910 -50210 2911 -47302
rect -3011 -50211 2911 -50210
rect -102 -50589 2 -50211
rect -3011 -50590 2911 -50589
rect -3011 -53498 -3010 -50590
rect -3200 -53602 -3010 -53498
rect -3011 -56510 -3010 -53602
rect 2910 -53498 2911 -50590
rect 2910 -53602 3100 -53498
rect 2910 -56510 2911 -53602
rect -3011 -56511 2911 -56510
rect -102 -56889 2 -56511
rect -3011 -56890 2911 -56889
rect -3011 -59798 -3010 -56890
rect -3200 -59902 -3010 -59798
rect -3011 -62810 -3010 -59902
rect 2910 -59798 2911 -56890
rect 2910 -59902 3100 -59798
rect 2910 -62810 2911 -59902
rect -3011 -62811 2911 -62810
rect -102 -63189 2 -62811
rect -3011 -63190 2911 -63189
rect -3011 -66098 -3010 -63190
rect -3200 -66202 -3010 -66098
rect -3011 -69110 -3010 -66202
rect 2910 -66098 2911 -63190
rect 2910 -66202 3100 -66098
rect 2910 -69110 2911 -66202
rect -3011 -69111 2911 -69110
rect -102 -69489 2 -69111
rect -3011 -69490 2911 -69489
rect -3011 -72398 -3010 -69490
rect -3200 -72502 -3010 -72398
rect -3011 -75410 -3010 -72502
rect 2910 -72398 2911 -69490
rect 2910 -72502 3100 -72398
rect 2910 -75410 2911 -72502
rect -3011 -75411 2911 -75410
rect -102 -75789 2 -75411
rect -3011 -75790 2911 -75789
rect -3011 -78698 -3010 -75790
rect -3200 -78802 -3010 -78698
rect -3011 -81710 -3010 -78802
rect 2910 -78698 2911 -75790
rect 2910 -78802 3100 -78698
rect 2910 -81710 2911 -78802
rect -3011 -81711 2911 -81710
rect -102 -82089 2 -81711
rect -3011 -82090 2911 -82089
rect -3011 -84998 -3010 -82090
rect -3200 -85102 -3010 -84998
rect -3011 -88010 -3010 -85102
rect 2910 -84998 2911 -82090
rect 2910 -85102 3100 -84998
rect 2910 -88010 2911 -85102
rect -3011 -88011 2911 -88010
rect -102 -88389 2 -88011
rect -3011 -88390 2911 -88389
rect -3011 -91298 -3010 -88390
rect -3200 -91402 -3010 -91298
rect -3011 -94310 -3010 -91402
rect 2910 -91298 2911 -88390
rect 2910 -91402 3100 -91298
rect 2910 -94310 2911 -91402
rect -3011 -94311 2911 -94310
rect -102 -94689 2 -94311
rect -3011 -94690 2911 -94689
rect -3011 -97598 -3010 -94690
rect -3200 -97702 -3010 -97598
rect -3011 -100610 -3010 -97702
rect 2910 -97598 2911 -94690
rect 2910 -97702 3100 -97598
rect 2910 -100610 2911 -97702
rect -3011 -100611 2911 -100610
rect -102 -100800 2 -100611
<< properties >>
string FIXED_BBOX -3150 94550 3050 100750
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 32 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
