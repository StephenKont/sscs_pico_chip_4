magic
tech sky130A
magscale 1 2
timestamp 1665943203
<< error_p >>
rect -287 369 -225 375
rect -159 369 -97 375
rect -31 369 31 375
rect 97 369 159 375
rect 225 369 287 375
rect -287 335 -275 369
rect -159 335 -147 369
rect -31 335 -19 369
rect 97 335 109 369
rect 225 335 237 369
rect -287 329 -225 335
rect -159 329 -97 335
rect -31 329 31 335
rect 97 329 159 335
rect 225 329 287 335
rect -287 -335 -225 -329
rect -159 -335 -97 -329
rect -31 -335 31 -329
rect 97 -335 159 -329
rect 225 -335 287 -329
rect -287 -369 -275 -335
rect -159 -369 -147 -335
rect -31 -369 -19 -335
rect 97 -369 109 -335
rect 225 -369 237 -335
rect -287 -375 -225 -369
rect -159 -375 -97 -369
rect -31 -375 31 -369
rect 97 -375 159 -369
rect 225 -375 287 -369
<< nwell >>
rect -487 -507 487 507
<< pmoslvt >>
rect -291 -288 -221 288
rect -163 -288 -93 288
rect -35 -288 35 288
rect 93 -288 163 288
rect 221 -288 291 288
<< pdiff >>
rect -349 276 -291 288
rect -349 -276 -337 276
rect -303 -276 -291 276
rect -349 -288 -291 -276
rect -221 276 -163 288
rect -221 -276 -209 276
rect -175 -276 -163 276
rect -221 -288 -163 -276
rect -93 276 -35 288
rect -93 -276 -81 276
rect -47 -276 -35 276
rect -93 -288 -35 -276
rect 35 276 93 288
rect 35 -276 47 276
rect 81 -276 93 276
rect 35 -288 93 -276
rect 163 276 221 288
rect 163 -276 175 276
rect 209 -276 221 276
rect 163 -288 221 -276
rect 291 276 349 288
rect 291 -276 303 276
rect 337 -276 349 276
rect 291 -288 349 -276
<< pdiffc >>
rect -337 -276 -303 276
rect -209 -276 -175 276
rect -81 -276 -47 276
rect 47 -276 81 276
rect 175 -276 209 276
rect 303 -276 337 276
<< nsubdiff >>
rect -451 437 -355 471
rect 355 437 451 471
rect -451 375 -417 437
rect 417 375 451 437
rect -451 -437 -417 -375
rect 417 -437 451 -375
rect -451 -471 -355 -437
rect 355 -471 451 -437
<< nsubdiffcont >>
rect -355 437 355 471
rect -451 -375 -417 375
rect 417 -375 451 375
rect -355 -471 355 -437
<< poly >>
rect -291 369 -221 385
rect -291 335 -275 369
rect -237 335 -221 369
rect -291 288 -221 335
rect -163 369 -93 385
rect -163 335 -147 369
rect -109 335 -93 369
rect -163 288 -93 335
rect -35 369 35 385
rect -35 335 -19 369
rect 19 335 35 369
rect -35 288 35 335
rect 93 369 163 385
rect 93 335 109 369
rect 147 335 163 369
rect 93 288 163 335
rect 221 369 291 385
rect 221 335 237 369
rect 275 335 291 369
rect 221 288 291 335
rect -291 -335 -221 -288
rect -291 -369 -275 -335
rect -237 -369 -221 -335
rect -291 -385 -221 -369
rect -163 -335 -93 -288
rect -163 -369 -147 -335
rect -109 -369 -93 -335
rect -163 -385 -93 -369
rect -35 -335 35 -288
rect -35 -369 -19 -335
rect 19 -369 35 -335
rect -35 -385 35 -369
rect 93 -335 163 -288
rect 93 -369 109 -335
rect 147 -369 163 -335
rect 93 -385 163 -369
rect 221 -335 291 -288
rect 221 -369 237 -335
rect 275 -369 291 -335
rect 221 -385 291 -369
<< polycont >>
rect -275 335 -237 369
rect -147 335 -109 369
rect -19 335 19 369
rect 109 335 147 369
rect 237 335 275 369
rect -275 -369 -237 -335
rect -147 -369 -109 -335
rect -19 -369 19 -335
rect 109 -369 147 -335
rect 237 -369 275 -335
<< locali >>
rect -451 437 -355 471
rect 355 437 451 471
rect -451 375 -417 437
rect 417 375 451 437
rect -291 335 -275 369
rect -237 335 -221 369
rect -163 335 -147 369
rect -109 335 -93 369
rect -35 335 -19 369
rect 19 335 35 369
rect 93 335 109 369
rect 147 335 163 369
rect 221 335 237 369
rect 275 335 291 369
rect -337 276 -303 292
rect -337 -292 -303 -276
rect -209 276 -175 292
rect -209 -292 -175 -276
rect -81 276 -47 292
rect -81 -292 -47 -276
rect 47 276 81 292
rect 47 -292 81 -276
rect 175 276 209 292
rect 175 -292 209 -276
rect 303 276 337 292
rect 303 -292 337 -276
rect -291 -369 -275 -335
rect -237 -369 -221 -335
rect -163 -369 -147 -335
rect -109 -369 -93 -335
rect -35 -369 -19 -335
rect 19 -369 35 -335
rect 93 -369 109 -335
rect 147 -369 163 -335
rect 221 -369 237 -335
rect 275 -369 291 -335
rect -451 -437 -417 -375
rect 417 -437 451 -375
rect -451 -471 -355 -437
rect 355 -471 451 -437
<< viali >>
rect -275 335 -237 369
rect -147 335 -109 369
rect -19 335 19 369
rect 109 335 147 369
rect 237 335 275 369
rect -337 -276 -303 276
rect -209 -276 -175 276
rect -81 -276 -47 276
rect 47 -276 81 276
rect 175 -276 209 276
rect 303 -276 337 276
rect -275 -369 -237 -335
rect -147 -369 -109 -335
rect -19 -369 19 -335
rect 109 -369 147 -335
rect 237 -369 275 -335
<< metal1 >>
rect -287 369 -225 375
rect -287 335 -275 369
rect -237 335 -225 369
rect -287 329 -225 335
rect -159 369 -97 375
rect -159 335 -147 369
rect -109 335 -97 369
rect -159 329 -97 335
rect -31 369 31 375
rect -31 335 -19 369
rect 19 335 31 369
rect -31 329 31 335
rect 97 369 159 375
rect 97 335 109 369
rect 147 335 159 369
rect 97 329 159 335
rect 225 369 287 375
rect 225 335 237 369
rect 275 335 287 369
rect 225 329 287 335
rect -343 276 -297 288
rect -343 -276 -337 276
rect -303 -276 -297 276
rect -343 -288 -297 -276
rect -215 276 -169 288
rect -215 -276 -209 276
rect -175 -276 -169 276
rect -215 -288 -169 -276
rect -87 276 -41 288
rect -87 -276 -81 276
rect -47 -276 -41 276
rect -87 -288 -41 -276
rect 41 276 87 288
rect 41 -276 47 276
rect 81 -276 87 276
rect 41 -288 87 -276
rect 169 276 215 288
rect 169 -276 175 276
rect 209 -276 215 276
rect 169 -288 215 -276
rect 297 276 343 288
rect 297 -276 303 276
rect 337 -276 343 276
rect 297 -288 343 -276
rect -287 -335 -225 -329
rect -287 -369 -275 -335
rect -237 -369 -225 -335
rect -287 -375 -225 -369
rect -159 -335 -97 -329
rect -159 -369 -147 -335
rect -109 -369 -97 -335
rect -159 -375 -97 -369
rect -31 -335 31 -329
rect -31 -369 -19 -335
rect 19 -369 31 -335
rect -31 -375 31 -369
rect 97 -335 159 -329
rect 97 -369 109 -335
rect 147 -369 159 -335
rect 97 -375 159 -369
rect 225 -335 287 -329
rect 225 -369 237 -335
rect 275 -369 287 -335
rect 225 -375 287 -369
<< properties >>
string FIXED_BBOX -434 -454 434 454
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2.88 l 0.35 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
