magic
tech sky130A
magscale 1 2
timestamp 1668293870
<< pwell >>
rect -321 -710 321 710
<< nmos >>
rect -125 -500 125 500
<< ndiff >>
rect -183 488 -125 500
rect -183 -488 -171 488
rect -137 -488 -125 488
rect -183 -500 -125 -488
rect 125 488 183 500
rect 125 -488 137 488
rect 171 -488 183 488
rect 125 -500 183 -488
<< ndiffc >>
rect -171 -488 -137 488
rect 137 -488 171 488
<< psubdiff >>
rect -285 640 -189 674
rect 189 640 285 674
rect -285 578 -251 640
rect 251 578 285 640
rect -285 -640 -251 -578
rect 251 -640 285 -578
rect -285 -674 -189 -640
rect 189 -674 285 -640
<< psubdiffcont >>
rect -189 640 189 674
rect -285 -578 -251 578
rect 251 -578 285 578
rect -189 -674 189 -640
<< poly >>
rect -125 572 125 588
rect -125 538 -109 572
rect 109 538 125 572
rect -125 500 125 538
rect -125 -538 125 -500
rect -125 -572 -109 -538
rect 109 -572 125 -538
rect -125 -588 125 -572
<< polycont >>
rect -109 538 109 572
rect -109 -572 109 -538
<< locali >>
rect -285 640 -189 674
rect 189 640 285 674
rect -285 578 -251 640
rect 251 578 285 640
rect -125 538 -109 572
rect 109 538 125 572
rect -171 488 -137 504
rect -171 -504 -137 -488
rect 137 488 171 504
rect 137 -504 171 -488
rect -125 -572 -109 -538
rect 109 -572 125 -538
rect -285 -640 -251 -578
rect 251 -640 285 -578
rect -285 -674 -189 -640
rect 189 -674 285 -640
<< viali >>
rect -109 538 109 572
rect -171 -488 -137 488
rect 137 -488 171 488
rect -109 -572 109 -538
<< metal1 >>
rect -121 572 121 578
rect -121 538 -109 572
rect 109 538 121 572
rect -121 532 121 538
rect -177 488 -131 500
rect -177 -488 -171 488
rect -137 -488 -131 488
rect -177 -500 -131 -488
rect 131 488 177 500
rect 131 -488 137 488
rect 171 -488 177 488
rect 131 -500 177 -488
rect -121 -538 121 -532
rect -121 -572 -109 -538
rect 109 -572 121 -538
rect -121 -578 121 -572
<< properties >>
string FIXED_BBOX -268 -657 268 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 1.25 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
