magic
tech sky130A
magscale 1 2
timestamp 1665339416
<< metal4 >>
rect -1351 2059 1351 2100
rect -1351 -2059 1095 2059
rect 1331 -2059 1351 2059
rect -1351 -2100 1351 -2059
<< via4 >>
rect 1095 -2059 1331 2059
<< mimcap2 >>
rect -1251 1960 749 2000
rect -1251 -1960 -1211 1960
rect 709 -1960 749 1960
rect -1251 -2000 749 -1960
<< mimcap2contact >>
rect -1211 -1960 709 1960
<< metal5 >>
rect 1053 2059 1373 2101
rect -1235 1960 733 1984
rect -1235 -1960 -1211 1960
rect 709 -1960 733 1960
rect -1235 -1984 733 -1960
rect 1053 -2059 1095 2059
rect 1331 -2059 1373 2059
rect 1053 -2101 1373 -2059
<< properties >>
string FIXED_BBOX -1351 -2100 849 2100
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 10 l 20 val 411.4 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
