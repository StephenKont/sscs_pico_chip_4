magic
tech sky130A
timestamp 1665170787
<< nwell >>
rect -1396 -1396 1396 1396
<< pwell >>
rect -1486 1396 1486 1486
rect -1486 -1396 -1396 1396
rect 1396 -1396 1486 1396
rect -1486 -1486 1486 -1396
<< mvpsubdiff >>
rect -1468 1462 1468 1468
rect -1468 1445 -1414 1462
rect 1414 1445 1468 1462
rect -1468 1439 1468 1445
rect -1468 1414 -1439 1439
rect -1468 -1414 -1462 1414
rect -1445 -1414 -1439 1414
rect 1439 1414 1468 1439
rect -1468 -1439 -1439 -1414
rect 1439 -1414 1445 1414
rect 1462 -1414 1468 1414
rect 1439 -1439 1468 -1414
rect -1468 -1445 1468 -1439
rect -1468 -1462 -1414 -1445
rect 1414 -1462 1468 -1445
rect -1468 -1468 1468 -1462
<< mvnsubdiff >>
rect -1363 1357 -731 1363
rect -1363 1340 -1309 1357
rect -785 1340 -731 1357
rect -1363 1334 -731 1340
rect -1363 1309 -1334 1334
rect -1363 785 -1357 1309
rect -1340 785 -1334 1309
rect -760 1309 -731 1334
rect -1363 760 -1334 785
rect -760 785 -754 1309
rect -737 785 -731 1309
rect -760 760 -731 785
rect -1363 754 -731 760
rect -1363 737 -1309 754
rect -785 737 -731 754
rect -1363 731 -731 737
rect -665 1357 -33 1363
rect -665 1340 -611 1357
rect -87 1340 -33 1357
rect -665 1334 -33 1340
rect -665 1309 -636 1334
rect -665 785 -659 1309
rect -642 785 -636 1309
rect -62 1309 -33 1334
rect -665 760 -636 785
rect -62 785 -56 1309
rect -39 785 -33 1309
rect -62 760 -33 785
rect -665 754 -33 760
rect -665 737 -611 754
rect -87 737 -33 754
rect -665 731 -33 737
rect 33 1357 665 1363
rect 33 1340 87 1357
rect 611 1340 665 1357
rect 33 1334 665 1340
rect 33 1309 62 1334
rect 33 785 39 1309
rect 56 785 62 1309
rect 636 1309 665 1334
rect 33 760 62 785
rect 636 785 642 1309
rect 659 785 665 1309
rect 636 760 665 785
rect 33 754 665 760
rect 33 737 87 754
rect 611 737 665 754
rect 33 731 665 737
rect 731 1357 1363 1363
rect 731 1340 785 1357
rect 1309 1340 1363 1357
rect 731 1334 1363 1340
rect 731 1309 760 1334
rect 731 785 737 1309
rect 754 785 760 1309
rect 1334 1309 1363 1334
rect 731 760 760 785
rect 1334 785 1340 1309
rect 1357 785 1363 1309
rect 1334 760 1363 785
rect 731 754 1363 760
rect 731 737 785 754
rect 1309 737 1363 754
rect 731 731 1363 737
rect -1363 659 -731 665
rect -1363 642 -1309 659
rect -785 642 -731 659
rect -1363 636 -731 642
rect -1363 611 -1334 636
rect -1363 87 -1357 611
rect -1340 87 -1334 611
rect -760 611 -731 636
rect -1363 62 -1334 87
rect -760 87 -754 611
rect -737 87 -731 611
rect -760 62 -731 87
rect -1363 56 -731 62
rect -1363 39 -1309 56
rect -785 39 -731 56
rect -1363 33 -731 39
rect -665 659 -33 665
rect -665 642 -611 659
rect -87 642 -33 659
rect -665 636 -33 642
rect -665 611 -636 636
rect -665 87 -659 611
rect -642 87 -636 611
rect -62 611 -33 636
rect -665 62 -636 87
rect -62 87 -56 611
rect -39 87 -33 611
rect -62 62 -33 87
rect -665 56 -33 62
rect -665 39 -611 56
rect -87 39 -33 56
rect -665 33 -33 39
rect 33 659 665 665
rect 33 642 87 659
rect 611 642 665 659
rect 33 636 665 642
rect 33 611 62 636
rect 33 87 39 611
rect 56 87 62 611
rect 636 611 665 636
rect 33 62 62 87
rect 636 87 642 611
rect 659 87 665 611
rect 636 62 665 87
rect 33 56 665 62
rect 33 39 87 56
rect 611 39 665 56
rect 33 33 665 39
rect 731 659 1363 665
rect 731 642 785 659
rect 1309 642 1363 659
rect 731 636 1363 642
rect 731 611 760 636
rect 731 87 737 611
rect 754 87 760 611
rect 1334 611 1363 636
rect 731 62 760 87
rect 1334 87 1340 611
rect 1357 87 1363 611
rect 1334 62 1363 87
rect 731 56 1363 62
rect 731 39 785 56
rect 1309 39 1363 56
rect 731 33 1363 39
rect -1363 -39 -731 -33
rect -1363 -56 -1309 -39
rect -785 -56 -731 -39
rect -1363 -62 -731 -56
rect -1363 -87 -1334 -62
rect -1363 -611 -1357 -87
rect -1340 -611 -1334 -87
rect -760 -87 -731 -62
rect -1363 -636 -1334 -611
rect -760 -611 -754 -87
rect -737 -611 -731 -87
rect -760 -636 -731 -611
rect -1363 -642 -731 -636
rect -1363 -659 -1309 -642
rect -785 -659 -731 -642
rect -1363 -665 -731 -659
rect -665 -39 -33 -33
rect -665 -56 -611 -39
rect -87 -56 -33 -39
rect -665 -62 -33 -56
rect -665 -87 -636 -62
rect -665 -611 -659 -87
rect -642 -611 -636 -87
rect -62 -87 -33 -62
rect -665 -636 -636 -611
rect -62 -611 -56 -87
rect -39 -611 -33 -87
rect -62 -636 -33 -611
rect -665 -642 -33 -636
rect -665 -659 -611 -642
rect -87 -659 -33 -642
rect -665 -665 -33 -659
rect 33 -39 665 -33
rect 33 -56 87 -39
rect 611 -56 665 -39
rect 33 -62 665 -56
rect 33 -87 62 -62
rect 33 -611 39 -87
rect 56 -611 62 -87
rect 636 -87 665 -62
rect 33 -636 62 -611
rect 636 -611 642 -87
rect 659 -611 665 -87
rect 636 -636 665 -611
rect 33 -642 665 -636
rect 33 -659 87 -642
rect 611 -659 665 -642
rect 33 -665 665 -659
rect 731 -39 1363 -33
rect 731 -56 785 -39
rect 1309 -56 1363 -39
rect 731 -62 1363 -56
rect 731 -87 760 -62
rect 731 -611 737 -87
rect 754 -611 760 -87
rect 1334 -87 1363 -62
rect 731 -636 760 -611
rect 1334 -611 1340 -87
rect 1357 -611 1363 -87
rect 1334 -636 1363 -611
rect 731 -642 1363 -636
rect 731 -659 785 -642
rect 1309 -659 1363 -642
rect 731 -665 1363 -659
rect -1363 -737 -731 -731
rect -1363 -754 -1309 -737
rect -785 -754 -731 -737
rect -1363 -760 -731 -754
rect -1363 -785 -1334 -760
rect -1363 -1309 -1357 -785
rect -1340 -1309 -1334 -785
rect -760 -785 -731 -760
rect -1363 -1334 -1334 -1309
rect -760 -1309 -754 -785
rect -737 -1309 -731 -785
rect -760 -1334 -731 -1309
rect -1363 -1340 -731 -1334
rect -1363 -1357 -1309 -1340
rect -785 -1357 -731 -1340
rect -1363 -1363 -731 -1357
rect -665 -737 -33 -731
rect -665 -754 -611 -737
rect -87 -754 -33 -737
rect -665 -760 -33 -754
rect -665 -785 -636 -760
rect -665 -1309 -659 -785
rect -642 -1309 -636 -785
rect -62 -785 -33 -760
rect -665 -1334 -636 -1309
rect -62 -1309 -56 -785
rect -39 -1309 -33 -785
rect -62 -1334 -33 -1309
rect -665 -1340 -33 -1334
rect -665 -1357 -611 -1340
rect -87 -1357 -33 -1340
rect -665 -1363 -33 -1357
rect 33 -737 665 -731
rect 33 -754 87 -737
rect 611 -754 665 -737
rect 33 -760 665 -754
rect 33 -785 62 -760
rect 33 -1309 39 -785
rect 56 -1309 62 -785
rect 636 -785 665 -760
rect 33 -1334 62 -1309
rect 636 -1309 642 -785
rect 659 -1309 665 -785
rect 636 -1334 665 -1309
rect 33 -1340 665 -1334
rect 33 -1357 87 -1340
rect 611 -1357 665 -1340
rect 33 -1363 665 -1357
rect 731 -737 1363 -731
rect 731 -754 785 -737
rect 1309 -754 1363 -737
rect 731 -760 1363 -754
rect 731 -785 760 -760
rect 731 -1309 737 -785
rect 754 -1309 760 -785
rect 1334 -785 1363 -760
rect 731 -1334 760 -1309
rect 1334 -1309 1340 -785
rect 1357 -1309 1363 -785
rect 1334 -1334 1363 -1309
rect 731 -1340 1363 -1334
rect 731 -1357 785 -1340
rect 1309 -1357 1363 -1340
rect 731 -1363 1363 -1357
<< mvpsubdiffcont >>
rect -1414 1445 1414 1462
rect -1462 -1414 -1445 1414
rect 1445 -1414 1462 1414
rect -1414 -1462 1414 -1445
<< mvnsubdiffcont >>
rect -1309 1340 -785 1357
rect -1357 785 -1340 1309
rect -754 785 -737 1309
rect -1309 737 -785 754
rect -611 1340 -87 1357
rect -659 785 -642 1309
rect -56 785 -39 1309
rect -611 737 -87 754
rect 87 1340 611 1357
rect 39 785 56 1309
rect 642 785 659 1309
rect 87 737 611 754
rect 785 1340 1309 1357
rect 737 785 754 1309
rect 1340 785 1357 1309
rect 785 737 1309 754
rect -1309 642 -785 659
rect -1357 87 -1340 611
rect -754 87 -737 611
rect -1309 39 -785 56
rect -611 642 -87 659
rect -659 87 -642 611
rect -56 87 -39 611
rect -611 39 -87 56
rect 87 642 611 659
rect 39 87 56 611
rect 642 87 659 611
rect 87 39 611 56
rect 785 642 1309 659
rect 737 87 754 611
rect 1340 87 1357 611
rect 785 39 1309 56
rect -1309 -56 -785 -39
rect -1357 -611 -1340 -87
rect -754 -611 -737 -87
rect -1309 -659 -785 -642
rect -611 -56 -87 -39
rect -659 -611 -642 -87
rect -56 -611 -39 -87
rect -611 -659 -87 -642
rect 87 -56 611 -39
rect 39 -611 56 -87
rect 642 -611 659 -87
rect 87 -659 611 -642
rect 785 -56 1309 -39
rect 737 -611 754 -87
rect 1340 -611 1357 -87
rect 785 -659 1309 -642
rect -1309 -754 -785 -737
rect -1357 -1309 -1340 -785
rect -754 -1309 -737 -785
rect -1309 -1357 -785 -1340
rect -611 -754 -87 -737
rect -659 -1309 -642 -785
rect -56 -1309 -39 -785
rect -611 -1357 -87 -1340
rect 87 -754 611 -737
rect 39 -1309 56 -785
rect 642 -1309 659 -785
rect 87 -1357 611 -1340
rect 785 -754 1309 -737
rect 737 -1309 754 -785
rect 1340 -1309 1357 -785
rect 785 -1357 1309 -1340
<< mvpdiode >>
rect -1297 1291 -797 1297
rect -1297 803 -1291 1291
rect -803 803 -797 1291
rect -1297 797 -797 803
rect -599 1291 -99 1297
rect -599 803 -593 1291
rect -105 803 -99 1291
rect -599 797 -99 803
rect 99 1291 599 1297
rect 99 803 105 1291
rect 593 803 599 1291
rect 99 797 599 803
rect 797 1291 1297 1297
rect 797 803 803 1291
rect 1291 803 1297 1291
rect 797 797 1297 803
rect -1297 593 -797 599
rect -1297 105 -1291 593
rect -803 105 -797 593
rect -1297 99 -797 105
rect -599 593 -99 599
rect -599 105 -593 593
rect -105 105 -99 593
rect -599 99 -99 105
rect 99 593 599 599
rect 99 105 105 593
rect 593 105 599 593
rect 99 99 599 105
rect 797 593 1297 599
rect 797 105 803 593
rect 1291 105 1297 593
rect 797 99 1297 105
rect -1297 -105 -797 -99
rect -1297 -593 -1291 -105
rect -803 -593 -797 -105
rect -1297 -599 -797 -593
rect -599 -105 -99 -99
rect -599 -593 -593 -105
rect -105 -593 -99 -105
rect -599 -599 -99 -593
rect 99 -105 599 -99
rect 99 -593 105 -105
rect 593 -593 599 -105
rect 99 -599 599 -593
rect 797 -105 1297 -99
rect 797 -593 803 -105
rect 1291 -593 1297 -105
rect 797 -599 1297 -593
rect -1297 -803 -797 -797
rect -1297 -1291 -1291 -803
rect -803 -1291 -797 -803
rect -1297 -1297 -797 -1291
rect -599 -803 -99 -797
rect -599 -1291 -593 -803
rect -105 -1291 -99 -803
rect -599 -1297 -99 -1291
rect 99 -803 599 -797
rect 99 -1291 105 -803
rect 593 -1291 599 -803
rect 99 -1297 599 -1291
rect 797 -803 1297 -797
rect 797 -1291 803 -803
rect 1291 -1291 1297 -803
rect 797 -1297 1297 -1291
<< mvpdiodec >>
rect -1291 803 -803 1291
rect -593 803 -105 1291
rect 105 803 593 1291
rect 803 803 1291 1291
rect -1291 105 -803 593
rect -593 105 -105 593
rect 105 105 593 593
rect 803 105 1291 593
rect -1291 -593 -803 -105
rect -593 -593 -105 -105
rect 105 -593 593 -105
rect 803 -593 1291 -105
rect -1291 -1291 -803 -803
rect -593 -1291 -105 -803
rect 105 -1291 593 -803
rect 803 -1291 1291 -803
<< locali >>
rect -1462 1445 -1414 1462
rect 1414 1445 1462 1462
rect -1462 1414 -1445 1445
rect 1445 1414 1462 1445
rect -1357 1340 -1309 1357
rect -785 1340 -737 1357
rect -1357 1309 -1340 1340
rect -754 1309 -737 1340
rect -1299 803 -1291 1291
rect -803 803 -795 1291
rect -1357 754 -1340 785
rect -754 754 -737 785
rect -1357 737 -1309 754
rect -785 737 -737 754
rect -659 1340 -611 1357
rect -87 1340 -39 1357
rect -659 1309 -642 1340
rect -56 1309 -39 1340
rect -601 803 -593 1291
rect -105 803 -97 1291
rect -659 754 -642 785
rect -56 754 -39 785
rect -659 737 -611 754
rect -87 737 -39 754
rect 39 1340 87 1357
rect 611 1340 659 1357
rect 39 1309 56 1340
rect 642 1309 659 1340
rect 97 803 105 1291
rect 593 803 601 1291
rect 39 754 56 785
rect 642 754 659 785
rect 39 737 87 754
rect 611 737 659 754
rect 737 1340 785 1357
rect 1309 1340 1357 1357
rect 737 1309 754 1340
rect 1340 1309 1357 1340
rect 795 803 803 1291
rect 1291 803 1299 1291
rect 737 754 754 785
rect 1340 754 1357 785
rect 737 737 785 754
rect 1309 737 1357 754
rect -1357 642 -1309 659
rect -785 642 -737 659
rect -1357 611 -1340 642
rect -754 611 -737 642
rect -1299 105 -1291 593
rect -803 105 -795 593
rect -1357 56 -1340 87
rect -754 56 -737 87
rect -1357 39 -1309 56
rect -785 39 -737 56
rect -659 642 -611 659
rect -87 642 -39 659
rect -659 611 -642 642
rect -56 611 -39 642
rect -601 105 -593 593
rect -105 105 -97 593
rect -659 56 -642 87
rect -56 56 -39 87
rect -659 39 -611 56
rect -87 39 -39 56
rect 39 642 87 659
rect 611 642 659 659
rect 39 611 56 642
rect 642 611 659 642
rect 97 105 105 593
rect 593 105 601 593
rect 39 56 56 87
rect 642 56 659 87
rect 39 39 87 56
rect 611 39 659 56
rect 737 642 785 659
rect 1309 642 1357 659
rect 737 611 754 642
rect 1340 611 1357 642
rect 795 105 803 593
rect 1291 105 1299 593
rect 737 56 754 87
rect 1340 56 1357 87
rect 737 39 785 56
rect 1309 39 1357 56
rect -1357 -56 -1309 -39
rect -785 -56 -737 -39
rect -1357 -87 -1340 -56
rect -754 -87 -737 -56
rect -1299 -593 -1291 -105
rect -803 -593 -795 -105
rect -1357 -642 -1340 -611
rect -754 -642 -737 -611
rect -1357 -659 -1309 -642
rect -785 -659 -737 -642
rect -659 -56 -611 -39
rect -87 -56 -39 -39
rect -659 -87 -642 -56
rect -56 -87 -39 -56
rect -601 -593 -593 -105
rect -105 -593 -97 -105
rect -659 -642 -642 -611
rect -56 -642 -39 -611
rect -659 -659 -611 -642
rect -87 -659 -39 -642
rect 39 -56 87 -39
rect 611 -56 659 -39
rect 39 -87 56 -56
rect 642 -87 659 -56
rect 97 -593 105 -105
rect 593 -593 601 -105
rect 39 -642 56 -611
rect 642 -642 659 -611
rect 39 -659 87 -642
rect 611 -659 659 -642
rect 737 -56 785 -39
rect 1309 -56 1357 -39
rect 737 -87 754 -56
rect 1340 -87 1357 -56
rect 795 -593 803 -105
rect 1291 -593 1299 -105
rect 737 -642 754 -611
rect 1340 -642 1357 -611
rect 737 -659 785 -642
rect 1309 -659 1357 -642
rect -1357 -754 -1309 -737
rect -785 -754 -737 -737
rect -1357 -785 -1340 -754
rect -754 -785 -737 -754
rect -1299 -1291 -1291 -803
rect -803 -1291 -795 -803
rect -1357 -1340 -1340 -1309
rect -754 -1340 -737 -1309
rect -1357 -1357 -1309 -1340
rect -785 -1357 -737 -1340
rect -659 -754 -611 -737
rect -87 -754 -39 -737
rect -659 -785 -642 -754
rect -56 -785 -39 -754
rect -601 -1291 -593 -803
rect -105 -1291 -97 -803
rect -659 -1340 -642 -1309
rect -56 -1340 -39 -1309
rect -659 -1357 -611 -1340
rect -87 -1357 -39 -1340
rect 39 -754 87 -737
rect 611 -754 659 -737
rect 39 -785 56 -754
rect 642 -785 659 -754
rect 97 -1291 105 -803
rect 593 -1291 601 -803
rect 39 -1340 56 -1309
rect 642 -1340 659 -1309
rect 39 -1357 87 -1340
rect 611 -1357 659 -1340
rect 737 -754 785 -737
rect 1309 -754 1357 -737
rect 737 -785 754 -754
rect 1340 -785 1357 -754
rect 795 -1291 803 -803
rect 1291 -1291 1299 -803
rect 737 -1340 754 -1309
rect 1340 -1340 1357 -1309
rect 737 -1357 785 -1340
rect 1309 -1357 1357 -1340
rect -1462 -1445 -1445 -1414
rect 1445 -1445 1462 -1414
rect -1462 -1462 -1414 -1445
rect 1414 -1462 1462 -1445
<< viali >>
rect -1291 803 -803 1291
rect -593 803 -105 1291
rect 105 803 593 1291
rect 803 803 1291 1291
rect -1291 105 -803 593
rect -593 105 -105 593
rect 105 105 593 593
rect 803 105 1291 593
rect -1291 -593 -803 -105
rect -593 -593 -105 -105
rect 105 -593 593 -105
rect 803 -593 1291 -105
rect -1291 -1291 -803 -803
rect -593 -1291 -105 -803
rect 105 -1291 593 -803
rect 803 -1291 1291 -803
<< metal1 >>
rect -1297 1291 -797 1294
rect -1297 803 -1291 1291
rect -803 803 -797 1291
rect -1297 800 -797 803
rect -599 1291 -99 1294
rect -599 803 -593 1291
rect -105 803 -99 1291
rect -599 800 -99 803
rect 99 1291 599 1294
rect 99 803 105 1291
rect 593 803 599 1291
rect 99 800 599 803
rect 797 1291 1297 1294
rect 797 803 803 1291
rect 1291 803 1297 1291
rect 797 800 1297 803
rect -1297 593 -797 596
rect -1297 105 -1291 593
rect -803 105 -797 593
rect -1297 102 -797 105
rect -599 593 -99 596
rect -599 105 -593 593
rect -105 105 -99 593
rect -599 102 -99 105
rect 99 593 599 596
rect 99 105 105 593
rect 593 105 599 593
rect 99 102 599 105
rect 797 593 1297 596
rect 797 105 803 593
rect 1291 105 1297 593
rect 797 102 1297 105
rect -1297 -105 -797 -102
rect -1297 -593 -1291 -105
rect -803 -593 -797 -105
rect -1297 -596 -797 -593
rect -599 -105 -99 -102
rect -599 -593 -593 -105
rect -105 -593 -99 -105
rect -599 -596 -99 -593
rect 99 -105 599 -102
rect 99 -593 105 -105
rect 593 -593 599 -105
rect 99 -596 599 -593
rect 797 -105 1297 -102
rect 797 -593 803 -105
rect 1291 -593 1297 -105
rect 797 -596 1297 -593
rect -1297 -803 -797 -800
rect -1297 -1291 -1291 -803
rect -803 -1291 -797 -803
rect -1297 -1294 -797 -1291
rect -599 -803 -99 -800
rect -599 -1291 -593 -803
rect -105 -1291 -99 -803
rect -599 -1294 -99 -1291
rect 99 -803 599 -800
rect 99 -1291 105 -803
rect 593 -1291 599 -803
rect 99 -1294 599 -1291
rect 797 -803 1297 -800
rect 797 -1291 803 -803
rect 1291 -1291 1297 -803
rect 797 -1294 1297 -1291
<< properties >>
string FIXED_BBOX 745 745 1348 1348
string gencell sky130_fd_pr__diode_pd2nw_11v0
string library sky130
string parameters w 5 l 5 area 25.0 peri 20.0 nx 4 ny 4 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 0 compatible {sky130_fd_pr__diode_pd2nw_05v5 sky130_fd_pr__diode_pd2nw_05v5_lvt  sky130_fd_pr__diode_pd2nw_05v5_hvt sky130_fd_pr__diode_pd2nw_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
