magic
tech sky130A
timestamp 1667516559
<< metal1 >>
rect 13991 -4393 54991 -4001
rect 13991 -13484 14525 -4393
rect 19548 -4543 54991 -4393
rect 19548 -13429 47532 -4543
rect 54381 -13429 54991 -4543
rect 19548 -13484 54991 -13429
rect 13991 -14001 54991 -13484
<< via1 >>
rect 14525 -13484 19548 -4393
rect 47532 -13429 54381 -4543
<< metal2 >>
rect 13991 -4393 54991 -4001
rect 13991 -13484 14525 -4393
rect 19548 -4543 54991 -4393
rect 19548 -13429 47532 -4543
rect 54381 -13429 54991 -4543
rect 19548 -13484 54991 -13429
rect 13991 -14001 54991 -13484
<< via2 >>
rect 14525 -13484 19548 -4393
rect 47532 -13429 54381 -4543
<< metal3 >>
rect 21491 40499 120491 48499
rect 13991 -4393 19991 -4001
rect 13991 -13484 14525 -4393
rect 19548 -13484 19991 -4393
rect 13991 -14001 19991 -13484
rect 21491 -4315 29491 40499
rect 21491 -13681 21873 -4315
rect 29086 -13681 29491 -4315
rect 21491 -14001 29491 -13681
rect 29991 31999 111991 39999
rect 29991 -44501 37991 31999
rect 38491 23499 103491 31499
rect 38491 -36001 46491 23499
rect 46991 -4543 54991 -4001
rect 46991 -13429 47532 -4543
rect 54381 -13429 54991 -4543
rect 46991 -27501 54991 -13429
rect 95491 -27501 103491 23499
rect 46991 -35501 103491 -27501
rect 103991 -36001 111991 31999
rect 38491 -44001 111991 -36001
rect 112491 -44501 120491 40499
rect 29991 -52501 120491 -44501
<< via3 >>
rect 14525 -13484 19548 -4393
rect 21873 -13681 29086 -4315
<< metal4 >>
rect 29991 40499 120491 48499
rect 13991 -4393 19991 -4001
rect 13991 -13484 14525 -4393
rect 19548 -13484 19991 -4393
rect 13991 -14001 19991 -13484
rect 21491 -4315 29491 -4001
rect 21491 -13681 21873 -4315
rect 29086 -13681 29491 -4315
rect 21491 -44501 29491 -13681
rect 29991 -36001 37991 40499
rect 38491 31999 111991 39999
rect 38491 -27501 46491 31999
rect 46991 23499 103491 31499
rect 46991 9493 54991 23499
rect 46991 676 47594 9493
rect 54457 676 54991 9493
rect 46991 -1 54991 676
rect 95491 -27501 103491 23499
rect 38491 -35501 103491 -27501
rect 103991 -36001 111991 31999
rect 29991 -44001 111991 -36001
rect 112491 -44501 120491 40499
rect 21491 -52501 120491 -44501
<< via4 >>
rect 14525 -13484 19548 -4393
rect 47594 676 54457 9493
<< metal5 >>
rect 21491 40499 120491 48499
rect 21491 9999 29491 40499
rect 13991 -1 29491 9999
rect 29991 31999 111991 39999
rect 13991 -4393 19991 -4001
rect 13991 -13484 14525 -4393
rect 19548 -13484 19991 -4393
rect 13991 -14001 19991 -13484
rect 29991 -44501 37991 31999
rect 38491 23499 103491 31499
rect 38491 -36001 46491 23499
rect 46991 9493 54991 9999
rect 46991 676 47594 9493
rect 54457 676 54991 9493
rect 46991 -27501 54991 676
rect 95491 -27501 103491 23499
rect 46991 -35501 103491 -27501
rect 103991 -36001 111991 31999
rect 38491 -44001 111991 -36001
rect 112491 -44501 120491 40499
rect 29991 -52501 120491 -44501
<< end >>
