magic
tech sky130A
magscale 1 2
timestamp 1665560017
<< nwell >>
rect -358 -1289 358 1289
<< mvpmos >>
rect -100 592 100 992
rect -100 64 100 464
rect -100 -464 100 -64
rect -100 -992 100 -592
<< mvpdiff >>
rect -158 980 -100 992
rect -158 604 -146 980
rect -112 604 -100 980
rect -158 592 -100 604
rect 100 980 158 992
rect 100 604 112 980
rect 146 604 158 980
rect 100 592 158 604
rect -158 452 -100 464
rect -158 76 -146 452
rect -112 76 -100 452
rect -158 64 -100 76
rect 100 452 158 464
rect 100 76 112 452
rect 146 76 158 452
rect 100 64 158 76
rect -158 -76 -100 -64
rect -158 -452 -146 -76
rect -112 -452 -100 -76
rect -158 -464 -100 -452
rect 100 -76 158 -64
rect 100 -452 112 -76
rect 146 -452 158 -76
rect 100 -464 158 -452
rect -158 -604 -100 -592
rect -158 -980 -146 -604
rect -112 -980 -100 -604
rect -158 -992 -100 -980
rect 100 -604 158 -592
rect 100 -980 112 -604
rect 146 -980 158 -604
rect 100 -992 158 -980
<< mvpdiffc >>
rect -146 604 -112 980
rect 112 604 146 980
rect -146 76 -112 452
rect 112 76 146 452
rect -146 -452 -112 -76
rect 112 -452 146 -76
rect -146 -980 -112 -604
rect 112 -980 146 -604
<< mvnsubdiff >>
rect -292 1211 292 1223
rect -292 1177 -184 1211
rect 184 1177 292 1211
rect -292 1165 292 1177
rect -292 1115 -234 1165
rect -292 -1115 -280 1115
rect -246 -1115 -234 1115
rect 234 1115 292 1165
rect -292 -1165 -234 -1115
rect 234 -1115 246 1115
rect 280 -1115 292 1115
rect 234 -1165 292 -1115
rect -292 -1177 292 -1165
rect -292 -1211 -184 -1177
rect 184 -1211 292 -1177
rect -292 -1223 292 -1211
<< mvnsubdiffcont >>
rect -184 1177 184 1211
rect -280 -1115 -246 1115
rect 246 -1115 280 1115
rect -184 -1211 184 -1177
<< poly >>
rect -100 1073 100 1089
rect -100 1039 -84 1073
rect 84 1039 100 1073
rect -100 992 100 1039
rect -100 545 100 592
rect -100 511 -84 545
rect 84 511 100 545
rect -100 464 100 511
rect -100 17 100 64
rect -100 -17 -84 17
rect 84 -17 100 17
rect -100 -64 100 -17
rect -100 -511 100 -464
rect -100 -545 -84 -511
rect 84 -545 100 -511
rect -100 -592 100 -545
rect -100 -1039 100 -992
rect -100 -1073 -84 -1039
rect 84 -1073 100 -1039
rect -100 -1089 100 -1073
<< polycont >>
rect -84 1039 84 1073
rect -84 511 84 545
rect -84 -17 84 17
rect -84 -545 84 -511
rect -84 -1073 84 -1039
<< locali >>
rect -280 1177 -184 1211
rect 184 1177 280 1211
rect -280 1115 -246 1177
rect 246 1115 280 1177
rect -100 1039 -84 1073
rect 84 1039 100 1073
rect -146 980 -112 996
rect -146 588 -112 604
rect 112 980 146 996
rect 112 588 146 604
rect -100 511 -84 545
rect 84 511 100 545
rect -146 452 -112 468
rect -146 60 -112 76
rect 112 452 146 468
rect 112 60 146 76
rect -100 -17 -84 17
rect 84 -17 100 17
rect -146 -76 -112 -60
rect -146 -468 -112 -452
rect 112 -76 146 -60
rect 112 -468 146 -452
rect -100 -545 -84 -511
rect 84 -545 100 -511
rect -146 -604 -112 -588
rect -146 -996 -112 -980
rect 112 -604 146 -588
rect 112 -996 146 -980
rect -100 -1073 -84 -1039
rect 84 -1073 100 -1039
rect -280 -1177 -246 -1115
rect 246 -1177 280 -1115
rect -280 -1211 -184 -1177
rect 184 -1211 280 -1177
<< viali >>
rect -84 1039 84 1073
rect -146 604 -112 980
rect 112 604 146 980
rect -84 511 84 545
rect -146 76 -112 452
rect 112 76 146 452
rect -84 -17 84 17
rect -146 -452 -112 -76
rect 112 -452 146 -76
rect -84 -545 84 -511
rect -146 -980 -112 -604
rect 112 -980 146 -604
rect -84 -1073 84 -1039
<< metal1 >>
rect -96 1073 96 1079
rect -96 1039 -84 1073
rect 84 1039 96 1073
rect -96 1033 96 1039
rect -152 980 -106 992
rect -152 604 -146 980
rect -112 604 -106 980
rect -152 592 -106 604
rect 106 980 152 992
rect 106 604 112 980
rect 146 604 152 980
rect 106 592 152 604
rect -96 545 96 551
rect -96 511 -84 545
rect 84 511 96 545
rect -96 505 96 511
rect -152 452 -106 464
rect -152 76 -146 452
rect -112 76 -106 452
rect -152 64 -106 76
rect 106 452 152 464
rect 106 76 112 452
rect 146 76 152 452
rect 106 64 152 76
rect -96 17 96 23
rect -96 -17 -84 17
rect 84 -17 96 17
rect -96 -23 96 -17
rect -152 -76 -106 -64
rect -152 -452 -146 -76
rect -112 -452 -106 -76
rect -152 -464 -106 -452
rect 106 -76 152 -64
rect 106 -452 112 -76
rect 146 -452 152 -76
rect 106 -464 152 -452
rect -96 -511 96 -505
rect -96 -545 -84 -511
rect 84 -545 96 -511
rect -96 -551 96 -545
rect -152 -604 -106 -592
rect -152 -980 -146 -604
rect -112 -980 -106 -604
rect -152 -992 -106 -980
rect 106 -604 152 -592
rect 106 -980 112 -604
rect 146 -980 152 -604
rect 106 -992 152 -980
rect -96 -1039 96 -1033
rect -96 -1073 -84 -1039
rect 84 -1073 96 -1039
rect -96 -1079 96 -1073
<< properties >>
string FIXED_BBOX -263 -1194 263 1194
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 1 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
