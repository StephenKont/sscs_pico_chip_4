magic
tech sky130A
magscale 1 2
timestamp 1666639277
<< nwell >>
rect -6549 -697 6549 697
<< mvpmos >>
rect -6291 -400 -6191 400
rect -6133 -400 -6033 400
rect -5975 -400 -5875 400
rect -5817 -400 -5717 400
rect -5659 -400 -5559 400
rect -5501 -400 -5401 400
rect -5343 -400 -5243 400
rect -5185 -400 -5085 400
rect -5027 -400 -4927 400
rect -4869 -400 -4769 400
rect -4711 -400 -4611 400
rect -4553 -400 -4453 400
rect -4395 -400 -4295 400
rect -4237 -400 -4137 400
rect -4079 -400 -3979 400
rect -3921 -400 -3821 400
rect -3763 -400 -3663 400
rect -3605 -400 -3505 400
rect -3447 -400 -3347 400
rect -3289 -400 -3189 400
rect -3131 -400 -3031 400
rect -2973 -400 -2873 400
rect -2815 -400 -2715 400
rect -2657 -400 -2557 400
rect -2499 -400 -2399 400
rect -2341 -400 -2241 400
rect -2183 -400 -2083 400
rect -2025 -400 -1925 400
rect -1867 -400 -1767 400
rect -1709 -400 -1609 400
rect -1551 -400 -1451 400
rect -1393 -400 -1293 400
rect -1235 -400 -1135 400
rect -1077 -400 -977 400
rect -919 -400 -819 400
rect -761 -400 -661 400
rect -603 -400 -503 400
rect -445 -400 -345 400
rect -287 -400 -187 400
rect -129 -400 -29 400
rect 29 -400 129 400
rect 187 -400 287 400
rect 345 -400 445 400
rect 503 -400 603 400
rect 661 -400 761 400
rect 819 -400 919 400
rect 977 -400 1077 400
rect 1135 -400 1235 400
rect 1293 -400 1393 400
rect 1451 -400 1551 400
rect 1609 -400 1709 400
rect 1767 -400 1867 400
rect 1925 -400 2025 400
rect 2083 -400 2183 400
rect 2241 -400 2341 400
rect 2399 -400 2499 400
rect 2557 -400 2657 400
rect 2715 -400 2815 400
rect 2873 -400 2973 400
rect 3031 -400 3131 400
rect 3189 -400 3289 400
rect 3347 -400 3447 400
rect 3505 -400 3605 400
rect 3663 -400 3763 400
rect 3821 -400 3921 400
rect 3979 -400 4079 400
rect 4137 -400 4237 400
rect 4295 -400 4395 400
rect 4453 -400 4553 400
rect 4611 -400 4711 400
rect 4769 -400 4869 400
rect 4927 -400 5027 400
rect 5085 -400 5185 400
rect 5243 -400 5343 400
rect 5401 -400 5501 400
rect 5559 -400 5659 400
rect 5717 -400 5817 400
rect 5875 -400 5975 400
rect 6033 -400 6133 400
rect 6191 -400 6291 400
<< mvpdiff >>
rect -6349 388 -6291 400
rect -6349 -388 -6337 388
rect -6303 -388 -6291 388
rect -6349 -400 -6291 -388
rect -6191 388 -6133 400
rect -6191 -388 -6179 388
rect -6145 -388 -6133 388
rect -6191 -400 -6133 -388
rect -6033 388 -5975 400
rect -6033 -388 -6021 388
rect -5987 -388 -5975 388
rect -6033 -400 -5975 -388
rect -5875 388 -5817 400
rect -5875 -388 -5863 388
rect -5829 -388 -5817 388
rect -5875 -400 -5817 -388
rect -5717 388 -5659 400
rect -5717 -388 -5705 388
rect -5671 -388 -5659 388
rect -5717 -400 -5659 -388
rect -5559 388 -5501 400
rect -5559 -388 -5547 388
rect -5513 -388 -5501 388
rect -5559 -400 -5501 -388
rect -5401 388 -5343 400
rect -5401 -388 -5389 388
rect -5355 -388 -5343 388
rect -5401 -400 -5343 -388
rect -5243 388 -5185 400
rect -5243 -388 -5231 388
rect -5197 -388 -5185 388
rect -5243 -400 -5185 -388
rect -5085 388 -5027 400
rect -5085 -388 -5073 388
rect -5039 -388 -5027 388
rect -5085 -400 -5027 -388
rect -4927 388 -4869 400
rect -4927 -388 -4915 388
rect -4881 -388 -4869 388
rect -4927 -400 -4869 -388
rect -4769 388 -4711 400
rect -4769 -388 -4757 388
rect -4723 -388 -4711 388
rect -4769 -400 -4711 -388
rect -4611 388 -4553 400
rect -4611 -388 -4599 388
rect -4565 -388 -4553 388
rect -4611 -400 -4553 -388
rect -4453 388 -4395 400
rect -4453 -388 -4441 388
rect -4407 -388 -4395 388
rect -4453 -400 -4395 -388
rect -4295 388 -4237 400
rect -4295 -388 -4283 388
rect -4249 -388 -4237 388
rect -4295 -400 -4237 -388
rect -4137 388 -4079 400
rect -4137 -388 -4125 388
rect -4091 -388 -4079 388
rect -4137 -400 -4079 -388
rect -3979 388 -3921 400
rect -3979 -388 -3967 388
rect -3933 -388 -3921 388
rect -3979 -400 -3921 -388
rect -3821 388 -3763 400
rect -3821 -388 -3809 388
rect -3775 -388 -3763 388
rect -3821 -400 -3763 -388
rect -3663 388 -3605 400
rect -3663 -388 -3651 388
rect -3617 -388 -3605 388
rect -3663 -400 -3605 -388
rect -3505 388 -3447 400
rect -3505 -388 -3493 388
rect -3459 -388 -3447 388
rect -3505 -400 -3447 -388
rect -3347 388 -3289 400
rect -3347 -388 -3335 388
rect -3301 -388 -3289 388
rect -3347 -400 -3289 -388
rect -3189 388 -3131 400
rect -3189 -388 -3177 388
rect -3143 -388 -3131 388
rect -3189 -400 -3131 -388
rect -3031 388 -2973 400
rect -3031 -388 -3019 388
rect -2985 -388 -2973 388
rect -3031 -400 -2973 -388
rect -2873 388 -2815 400
rect -2873 -388 -2861 388
rect -2827 -388 -2815 388
rect -2873 -400 -2815 -388
rect -2715 388 -2657 400
rect -2715 -388 -2703 388
rect -2669 -388 -2657 388
rect -2715 -400 -2657 -388
rect -2557 388 -2499 400
rect -2557 -388 -2545 388
rect -2511 -388 -2499 388
rect -2557 -400 -2499 -388
rect -2399 388 -2341 400
rect -2399 -388 -2387 388
rect -2353 -388 -2341 388
rect -2399 -400 -2341 -388
rect -2241 388 -2183 400
rect -2241 -388 -2229 388
rect -2195 -388 -2183 388
rect -2241 -400 -2183 -388
rect -2083 388 -2025 400
rect -2083 -388 -2071 388
rect -2037 -388 -2025 388
rect -2083 -400 -2025 -388
rect -1925 388 -1867 400
rect -1925 -388 -1913 388
rect -1879 -388 -1867 388
rect -1925 -400 -1867 -388
rect -1767 388 -1709 400
rect -1767 -388 -1755 388
rect -1721 -388 -1709 388
rect -1767 -400 -1709 -388
rect -1609 388 -1551 400
rect -1609 -388 -1597 388
rect -1563 -388 -1551 388
rect -1609 -400 -1551 -388
rect -1451 388 -1393 400
rect -1451 -388 -1439 388
rect -1405 -388 -1393 388
rect -1451 -400 -1393 -388
rect -1293 388 -1235 400
rect -1293 -388 -1281 388
rect -1247 -388 -1235 388
rect -1293 -400 -1235 -388
rect -1135 388 -1077 400
rect -1135 -388 -1123 388
rect -1089 -388 -1077 388
rect -1135 -400 -1077 -388
rect -977 388 -919 400
rect -977 -388 -965 388
rect -931 -388 -919 388
rect -977 -400 -919 -388
rect -819 388 -761 400
rect -819 -388 -807 388
rect -773 -388 -761 388
rect -819 -400 -761 -388
rect -661 388 -603 400
rect -661 -388 -649 388
rect -615 -388 -603 388
rect -661 -400 -603 -388
rect -503 388 -445 400
rect -503 -388 -491 388
rect -457 -388 -445 388
rect -503 -400 -445 -388
rect -345 388 -287 400
rect -345 -388 -333 388
rect -299 -388 -287 388
rect -345 -400 -287 -388
rect -187 388 -129 400
rect -187 -388 -175 388
rect -141 -388 -129 388
rect -187 -400 -129 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 129 388 187 400
rect 129 -388 141 388
rect 175 -388 187 388
rect 129 -400 187 -388
rect 287 388 345 400
rect 287 -388 299 388
rect 333 -388 345 388
rect 287 -400 345 -388
rect 445 388 503 400
rect 445 -388 457 388
rect 491 -388 503 388
rect 445 -400 503 -388
rect 603 388 661 400
rect 603 -388 615 388
rect 649 -388 661 388
rect 603 -400 661 -388
rect 761 388 819 400
rect 761 -388 773 388
rect 807 -388 819 388
rect 761 -400 819 -388
rect 919 388 977 400
rect 919 -388 931 388
rect 965 -388 977 388
rect 919 -400 977 -388
rect 1077 388 1135 400
rect 1077 -388 1089 388
rect 1123 -388 1135 388
rect 1077 -400 1135 -388
rect 1235 388 1293 400
rect 1235 -388 1247 388
rect 1281 -388 1293 388
rect 1235 -400 1293 -388
rect 1393 388 1451 400
rect 1393 -388 1405 388
rect 1439 -388 1451 388
rect 1393 -400 1451 -388
rect 1551 388 1609 400
rect 1551 -388 1563 388
rect 1597 -388 1609 388
rect 1551 -400 1609 -388
rect 1709 388 1767 400
rect 1709 -388 1721 388
rect 1755 -388 1767 388
rect 1709 -400 1767 -388
rect 1867 388 1925 400
rect 1867 -388 1879 388
rect 1913 -388 1925 388
rect 1867 -400 1925 -388
rect 2025 388 2083 400
rect 2025 -388 2037 388
rect 2071 -388 2083 388
rect 2025 -400 2083 -388
rect 2183 388 2241 400
rect 2183 -388 2195 388
rect 2229 -388 2241 388
rect 2183 -400 2241 -388
rect 2341 388 2399 400
rect 2341 -388 2353 388
rect 2387 -388 2399 388
rect 2341 -400 2399 -388
rect 2499 388 2557 400
rect 2499 -388 2511 388
rect 2545 -388 2557 388
rect 2499 -400 2557 -388
rect 2657 388 2715 400
rect 2657 -388 2669 388
rect 2703 -388 2715 388
rect 2657 -400 2715 -388
rect 2815 388 2873 400
rect 2815 -388 2827 388
rect 2861 -388 2873 388
rect 2815 -400 2873 -388
rect 2973 388 3031 400
rect 2973 -388 2985 388
rect 3019 -388 3031 388
rect 2973 -400 3031 -388
rect 3131 388 3189 400
rect 3131 -388 3143 388
rect 3177 -388 3189 388
rect 3131 -400 3189 -388
rect 3289 388 3347 400
rect 3289 -388 3301 388
rect 3335 -388 3347 388
rect 3289 -400 3347 -388
rect 3447 388 3505 400
rect 3447 -388 3459 388
rect 3493 -388 3505 388
rect 3447 -400 3505 -388
rect 3605 388 3663 400
rect 3605 -388 3617 388
rect 3651 -388 3663 388
rect 3605 -400 3663 -388
rect 3763 388 3821 400
rect 3763 -388 3775 388
rect 3809 -388 3821 388
rect 3763 -400 3821 -388
rect 3921 388 3979 400
rect 3921 -388 3933 388
rect 3967 -388 3979 388
rect 3921 -400 3979 -388
rect 4079 388 4137 400
rect 4079 -388 4091 388
rect 4125 -388 4137 388
rect 4079 -400 4137 -388
rect 4237 388 4295 400
rect 4237 -388 4249 388
rect 4283 -388 4295 388
rect 4237 -400 4295 -388
rect 4395 388 4453 400
rect 4395 -388 4407 388
rect 4441 -388 4453 388
rect 4395 -400 4453 -388
rect 4553 388 4611 400
rect 4553 -388 4565 388
rect 4599 -388 4611 388
rect 4553 -400 4611 -388
rect 4711 388 4769 400
rect 4711 -388 4723 388
rect 4757 -388 4769 388
rect 4711 -400 4769 -388
rect 4869 388 4927 400
rect 4869 -388 4881 388
rect 4915 -388 4927 388
rect 4869 -400 4927 -388
rect 5027 388 5085 400
rect 5027 -388 5039 388
rect 5073 -388 5085 388
rect 5027 -400 5085 -388
rect 5185 388 5243 400
rect 5185 -388 5197 388
rect 5231 -388 5243 388
rect 5185 -400 5243 -388
rect 5343 388 5401 400
rect 5343 -388 5355 388
rect 5389 -388 5401 388
rect 5343 -400 5401 -388
rect 5501 388 5559 400
rect 5501 -388 5513 388
rect 5547 -388 5559 388
rect 5501 -400 5559 -388
rect 5659 388 5717 400
rect 5659 -388 5671 388
rect 5705 -388 5717 388
rect 5659 -400 5717 -388
rect 5817 388 5875 400
rect 5817 -388 5829 388
rect 5863 -388 5875 388
rect 5817 -400 5875 -388
rect 5975 388 6033 400
rect 5975 -388 5987 388
rect 6021 -388 6033 388
rect 5975 -400 6033 -388
rect 6133 388 6191 400
rect 6133 -388 6145 388
rect 6179 -388 6191 388
rect 6133 -400 6191 -388
rect 6291 388 6349 400
rect 6291 -388 6303 388
rect 6337 -388 6349 388
rect 6291 -400 6349 -388
<< mvpdiffc >>
rect -6337 -388 -6303 388
rect -6179 -388 -6145 388
rect -6021 -388 -5987 388
rect -5863 -388 -5829 388
rect -5705 -388 -5671 388
rect -5547 -388 -5513 388
rect -5389 -388 -5355 388
rect -5231 -388 -5197 388
rect -5073 -388 -5039 388
rect -4915 -388 -4881 388
rect -4757 -388 -4723 388
rect -4599 -388 -4565 388
rect -4441 -388 -4407 388
rect -4283 -388 -4249 388
rect -4125 -388 -4091 388
rect -3967 -388 -3933 388
rect -3809 -388 -3775 388
rect -3651 -388 -3617 388
rect -3493 -388 -3459 388
rect -3335 -388 -3301 388
rect -3177 -388 -3143 388
rect -3019 -388 -2985 388
rect -2861 -388 -2827 388
rect -2703 -388 -2669 388
rect -2545 -388 -2511 388
rect -2387 -388 -2353 388
rect -2229 -388 -2195 388
rect -2071 -388 -2037 388
rect -1913 -388 -1879 388
rect -1755 -388 -1721 388
rect -1597 -388 -1563 388
rect -1439 -388 -1405 388
rect -1281 -388 -1247 388
rect -1123 -388 -1089 388
rect -965 -388 -931 388
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
rect 931 -388 965 388
rect 1089 -388 1123 388
rect 1247 -388 1281 388
rect 1405 -388 1439 388
rect 1563 -388 1597 388
rect 1721 -388 1755 388
rect 1879 -388 1913 388
rect 2037 -388 2071 388
rect 2195 -388 2229 388
rect 2353 -388 2387 388
rect 2511 -388 2545 388
rect 2669 -388 2703 388
rect 2827 -388 2861 388
rect 2985 -388 3019 388
rect 3143 -388 3177 388
rect 3301 -388 3335 388
rect 3459 -388 3493 388
rect 3617 -388 3651 388
rect 3775 -388 3809 388
rect 3933 -388 3967 388
rect 4091 -388 4125 388
rect 4249 -388 4283 388
rect 4407 -388 4441 388
rect 4565 -388 4599 388
rect 4723 -388 4757 388
rect 4881 -388 4915 388
rect 5039 -388 5073 388
rect 5197 -388 5231 388
rect 5355 -388 5389 388
rect 5513 -388 5547 388
rect 5671 -388 5705 388
rect 5829 -388 5863 388
rect 5987 -388 6021 388
rect 6145 -388 6179 388
rect 6303 -388 6337 388
<< mvnsubdiff >>
rect -6483 619 6483 631
rect -6483 585 -6375 619
rect 6375 585 6483 619
rect -6483 573 6483 585
rect -6483 523 -6425 573
rect -6483 -523 -6471 523
rect -6437 -523 -6425 523
rect 6425 523 6483 573
rect -6483 -573 -6425 -523
rect 6425 -523 6437 523
rect 6471 -523 6483 523
rect 6425 -573 6483 -523
rect -6483 -585 6483 -573
rect -6483 -619 -6375 -585
rect 6375 -619 6483 -585
rect -6483 -631 6483 -619
<< mvnsubdiffcont >>
rect -6375 585 6375 619
rect -6471 -523 -6437 523
rect 6437 -523 6471 523
rect -6375 -619 6375 -585
<< poly >>
rect -6291 481 -6191 497
rect -6291 447 -6275 481
rect -6207 447 -6191 481
rect -6291 400 -6191 447
rect -6133 481 -6033 497
rect -6133 447 -6117 481
rect -6049 447 -6033 481
rect -6133 400 -6033 447
rect -5975 481 -5875 497
rect -5975 447 -5959 481
rect -5891 447 -5875 481
rect -5975 400 -5875 447
rect -5817 481 -5717 497
rect -5817 447 -5801 481
rect -5733 447 -5717 481
rect -5817 400 -5717 447
rect -5659 481 -5559 497
rect -5659 447 -5643 481
rect -5575 447 -5559 481
rect -5659 400 -5559 447
rect -5501 481 -5401 497
rect -5501 447 -5485 481
rect -5417 447 -5401 481
rect -5501 400 -5401 447
rect -5343 481 -5243 497
rect -5343 447 -5327 481
rect -5259 447 -5243 481
rect -5343 400 -5243 447
rect -5185 481 -5085 497
rect -5185 447 -5169 481
rect -5101 447 -5085 481
rect -5185 400 -5085 447
rect -5027 481 -4927 497
rect -5027 447 -5011 481
rect -4943 447 -4927 481
rect -5027 400 -4927 447
rect -4869 481 -4769 497
rect -4869 447 -4853 481
rect -4785 447 -4769 481
rect -4869 400 -4769 447
rect -4711 481 -4611 497
rect -4711 447 -4695 481
rect -4627 447 -4611 481
rect -4711 400 -4611 447
rect -4553 481 -4453 497
rect -4553 447 -4537 481
rect -4469 447 -4453 481
rect -4553 400 -4453 447
rect -4395 481 -4295 497
rect -4395 447 -4379 481
rect -4311 447 -4295 481
rect -4395 400 -4295 447
rect -4237 481 -4137 497
rect -4237 447 -4221 481
rect -4153 447 -4137 481
rect -4237 400 -4137 447
rect -4079 481 -3979 497
rect -4079 447 -4063 481
rect -3995 447 -3979 481
rect -4079 400 -3979 447
rect -3921 481 -3821 497
rect -3921 447 -3905 481
rect -3837 447 -3821 481
rect -3921 400 -3821 447
rect -3763 481 -3663 497
rect -3763 447 -3747 481
rect -3679 447 -3663 481
rect -3763 400 -3663 447
rect -3605 481 -3505 497
rect -3605 447 -3589 481
rect -3521 447 -3505 481
rect -3605 400 -3505 447
rect -3447 481 -3347 497
rect -3447 447 -3431 481
rect -3363 447 -3347 481
rect -3447 400 -3347 447
rect -3289 481 -3189 497
rect -3289 447 -3273 481
rect -3205 447 -3189 481
rect -3289 400 -3189 447
rect -3131 481 -3031 497
rect -3131 447 -3115 481
rect -3047 447 -3031 481
rect -3131 400 -3031 447
rect -2973 481 -2873 497
rect -2973 447 -2957 481
rect -2889 447 -2873 481
rect -2973 400 -2873 447
rect -2815 481 -2715 497
rect -2815 447 -2799 481
rect -2731 447 -2715 481
rect -2815 400 -2715 447
rect -2657 481 -2557 497
rect -2657 447 -2641 481
rect -2573 447 -2557 481
rect -2657 400 -2557 447
rect -2499 481 -2399 497
rect -2499 447 -2483 481
rect -2415 447 -2399 481
rect -2499 400 -2399 447
rect -2341 481 -2241 497
rect -2341 447 -2325 481
rect -2257 447 -2241 481
rect -2341 400 -2241 447
rect -2183 481 -2083 497
rect -2183 447 -2167 481
rect -2099 447 -2083 481
rect -2183 400 -2083 447
rect -2025 481 -1925 497
rect -2025 447 -2009 481
rect -1941 447 -1925 481
rect -2025 400 -1925 447
rect -1867 481 -1767 497
rect -1867 447 -1851 481
rect -1783 447 -1767 481
rect -1867 400 -1767 447
rect -1709 481 -1609 497
rect -1709 447 -1693 481
rect -1625 447 -1609 481
rect -1709 400 -1609 447
rect -1551 481 -1451 497
rect -1551 447 -1535 481
rect -1467 447 -1451 481
rect -1551 400 -1451 447
rect -1393 481 -1293 497
rect -1393 447 -1377 481
rect -1309 447 -1293 481
rect -1393 400 -1293 447
rect -1235 481 -1135 497
rect -1235 447 -1219 481
rect -1151 447 -1135 481
rect -1235 400 -1135 447
rect -1077 481 -977 497
rect -1077 447 -1061 481
rect -993 447 -977 481
rect -1077 400 -977 447
rect -919 481 -819 497
rect -919 447 -903 481
rect -835 447 -819 481
rect -919 400 -819 447
rect -761 481 -661 497
rect -761 447 -745 481
rect -677 447 -661 481
rect -761 400 -661 447
rect -603 481 -503 497
rect -603 447 -587 481
rect -519 447 -503 481
rect -603 400 -503 447
rect -445 481 -345 497
rect -445 447 -429 481
rect -361 447 -345 481
rect -445 400 -345 447
rect -287 481 -187 497
rect -287 447 -271 481
rect -203 447 -187 481
rect -287 400 -187 447
rect -129 481 -29 497
rect -129 447 -113 481
rect -45 447 -29 481
rect -129 400 -29 447
rect 29 481 129 497
rect 29 447 45 481
rect 113 447 129 481
rect 29 400 129 447
rect 187 481 287 497
rect 187 447 203 481
rect 271 447 287 481
rect 187 400 287 447
rect 345 481 445 497
rect 345 447 361 481
rect 429 447 445 481
rect 345 400 445 447
rect 503 481 603 497
rect 503 447 519 481
rect 587 447 603 481
rect 503 400 603 447
rect 661 481 761 497
rect 661 447 677 481
rect 745 447 761 481
rect 661 400 761 447
rect 819 481 919 497
rect 819 447 835 481
rect 903 447 919 481
rect 819 400 919 447
rect 977 481 1077 497
rect 977 447 993 481
rect 1061 447 1077 481
rect 977 400 1077 447
rect 1135 481 1235 497
rect 1135 447 1151 481
rect 1219 447 1235 481
rect 1135 400 1235 447
rect 1293 481 1393 497
rect 1293 447 1309 481
rect 1377 447 1393 481
rect 1293 400 1393 447
rect 1451 481 1551 497
rect 1451 447 1467 481
rect 1535 447 1551 481
rect 1451 400 1551 447
rect 1609 481 1709 497
rect 1609 447 1625 481
rect 1693 447 1709 481
rect 1609 400 1709 447
rect 1767 481 1867 497
rect 1767 447 1783 481
rect 1851 447 1867 481
rect 1767 400 1867 447
rect 1925 481 2025 497
rect 1925 447 1941 481
rect 2009 447 2025 481
rect 1925 400 2025 447
rect 2083 481 2183 497
rect 2083 447 2099 481
rect 2167 447 2183 481
rect 2083 400 2183 447
rect 2241 481 2341 497
rect 2241 447 2257 481
rect 2325 447 2341 481
rect 2241 400 2341 447
rect 2399 481 2499 497
rect 2399 447 2415 481
rect 2483 447 2499 481
rect 2399 400 2499 447
rect 2557 481 2657 497
rect 2557 447 2573 481
rect 2641 447 2657 481
rect 2557 400 2657 447
rect 2715 481 2815 497
rect 2715 447 2731 481
rect 2799 447 2815 481
rect 2715 400 2815 447
rect 2873 481 2973 497
rect 2873 447 2889 481
rect 2957 447 2973 481
rect 2873 400 2973 447
rect 3031 481 3131 497
rect 3031 447 3047 481
rect 3115 447 3131 481
rect 3031 400 3131 447
rect 3189 481 3289 497
rect 3189 447 3205 481
rect 3273 447 3289 481
rect 3189 400 3289 447
rect 3347 481 3447 497
rect 3347 447 3363 481
rect 3431 447 3447 481
rect 3347 400 3447 447
rect 3505 481 3605 497
rect 3505 447 3521 481
rect 3589 447 3605 481
rect 3505 400 3605 447
rect 3663 481 3763 497
rect 3663 447 3679 481
rect 3747 447 3763 481
rect 3663 400 3763 447
rect 3821 481 3921 497
rect 3821 447 3837 481
rect 3905 447 3921 481
rect 3821 400 3921 447
rect 3979 481 4079 497
rect 3979 447 3995 481
rect 4063 447 4079 481
rect 3979 400 4079 447
rect 4137 481 4237 497
rect 4137 447 4153 481
rect 4221 447 4237 481
rect 4137 400 4237 447
rect 4295 481 4395 497
rect 4295 447 4311 481
rect 4379 447 4395 481
rect 4295 400 4395 447
rect 4453 481 4553 497
rect 4453 447 4469 481
rect 4537 447 4553 481
rect 4453 400 4553 447
rect 4611 481 4711 497
rect 4611 447 4627 481
rect 4695 447 4711 481
rect 4611 400 4711 447
rect 4769 481 4869 497
rect 4769 447 4785 481
rect 4853 447 4869 481
rect 4769 400 4869 447
rect 4927 481 5027 497
rect 4927 447 4943 481
rect 5011 447 5027 481
rect 4927 400 5027 447
rect 5085 481 5185 497
rect 5085 447 5101 481
rect 5169 447 5185 481
rect 5085 400 5185 447
rect 5243 481 5343 497
rect 5243 447 5259 481
rect 5327 447 5343 481
rect 5243 400 5343 447
rect 5401 481 5501 497
rect 5401 447 5417 481
rect 5485 447 5501 481
rect 5401 400 5501 447
rect 5559 481 5659 497
rect 5559 447 5575 481
rect 5643 447 5659 481
rect 5559 400 5659 447
rect 5717 481 5817 497
rect 5717 447 5733 481
rect 5801 447 5817 481
rect 5717 400 5817 447
rect 5875 481 5975 497
rect 5875 447 5891 481
rect 5959 447 5975 481
rect 5875 400 5975 447
rect 6033 481 6133 497
rect 6033 447 6049 481
rect 6117 447 6133 481
rect 6033 400 6133 447
rect 6191 481 6291 497
rect 6191 447 6207 481
rect 6275 447 6291 481
rect 6191 400 6291 447
rect -6291 -447 -6191 -400
rect -6291 -481 -6275 -447
rect -6207 -481 -6191 -447
rect -6291 -497 -6191 -481
rect -6133 -447 -6033 -400
rect -6133 -481 -6117 -447
rect -6049 -481 -6033 -447
rect -6133 -497 -6033 -481
rect -5975 -447 -5875 -400
rect -5975 -481 -5959 -447
rect -5891 -481 -5875 -447
rect -5975 -497 -5875 -481
rect -5817 -447 -5717 -400
rect -5817 -481 -5801 -447
rect -5733 -481 -5717 -447
rect -5817 -497 -5717 -481
rect -5659 -447 -5559 -400
rect -5659 -481 -5643 -447
rect -5575 -481 -5559 -447
rect -5659 -497 -5559 -481
rect -5501 -447 -5401 -400
rect -5501 -481 -5485 -447
rect -5417 -481 -5401 -447
rect -5501 -497 -5401 -481
rect -5343 -447 -5243 -400
rect -5343 -481 -5327 -447
rect -5259 -481 -5243 -447
rect -5343 -497 -5243 -481
rect -5185 -447 -5085 -400
rect -5185 -481 -5169 -447
rect -5101 -481 -5085 -447
rect -5185 -497 -5085 -481
rect -5027 -447 -4927 -400
rect -5027 -481 -5011 -447
rect -4943 -481 -4927 -447
rect -5027 -497 -4927 -481
rect -4869 -447 -4769 -400
rect -4869 -481 -4853 -447
rect -4785 -481 -4769 -447
rect -4869 -497 -4769 -481
rect -4711 -447 -4611 -400
rect -4711 -481 -4695 -447
rect -4627 -481 -4611 -447
rect -4711 -497 -4611 -481
rect -4553 -447 -4453 -400
rect -4553 -481 -4537 -447
rect -4469 -481 -4453 -447
rect -4553 -497 -4453 -481
rect -4395 -447 -4295 -400
rect -4395 -481 -4379 -447
rect -4311 -481 -4295 -447
rect -4395 -497 -4295 -481
rect -4237 -447 -4137 -400
rect -4237 -481 -4221 -447
rect -4153 -481 -4137 -447
rect -4237 -497 -4137 -481
rect -4079 -447 -3979 -400
rect -4079 -481 -4063 -447
rect -3995 -481 -3979 -447
rect -4079 -497 -3979 -481
rect -3921 -447 -3821 -400
rect -3921 -481 -3905 -447
rect -3837 -481 -3821 -447
rect -3921 -497 -3821 -481
rect -3763 -447 -3663 -400
rect -3763 -481 -3747 -447
rect -3679 -481 -3663 -447
rect -3763 -497 -3663 -481
rect -3605 -447 -3505 -400
rect -3605 -481 -3589 -447
rect -3521 -481 -3505 -447
rect -3605 -497 -3505 -481
rect -3447 -447 -3347 -400
rect -3447 -481 -3431 -447
rect -3363 -481 -3347 -447
rect -3447 -497 -3347 -481
rect -3289 -447 -3189 -400
rect -3289 -481 -3273 -447
rect -3205 -481 -3189 -447
rect -3289 -497 -3189 -481
rect -3131 -447 -3031 -400
rect -3131 -481 -3115 -447
rect -3047 -481 -3031 -447
rect -3131 -497 -3031 -481
rect -2973 -447 -2873 -400
rect -2973 -481 -2957 -447
rect -2889 -481 -2873 -447
rect -2973 -497 -2873 -481
rect -2815 -447 -2715 -400
rect -2815 -481 -2799 -447
rect -2731 -481 -2715 -447
rect -2815 -497 -2715 -481
rect -2657 -447 -2557 -400
rect -2657 -481 -2641 -447
rect -2573 -481 -2557 -447
rect -2657 -497 -2557 -481
rect -2499 -447 -2399 -400
rect -2499 -481 -2483 -447
rect -2415 -481 -2399 -447
rect -2499 -497 -2399 -481
rect -2341 -447 -2241 -400
rect -2341 -481 -2325 -447
rect -2257 -481 -2241 -447
rect -2341 -497 -2241 -481
rect -2183 -447 -2083 -400
rect -2183 -481 -2167 -447
rect -2099 -481 -2083 -447
rect -2183 -497 -2083 -481
rect -2025 -447 -1925 -400
rect -2025 -481 -2009 -447
rect -1941 -481 -1925 -447
rect -2025 -497 -1925 -481
rect -1867 -447 -1767 -400
rect -1867 -481 -1851 -447
rect -1783 -481 -1767 -447
rect -1867 -497 -1767 -481
rect -1709 -447 -1609 -400
rect -1709 -481 -1693 -447
rect -1625 -481 -1609 -447
rect -1709 -497 -1609 -481
rect -1551 -447 -1451 -400
rect -1551 -481 -1535 -447
rect -1467 -481 -1451 -447
rect -1551 -497 -1451 -481
rect -1393 -447 -1293 -400
rect -1393 -481 -1377 -447
rect -1309 -481 -1293 -447
rect -1393 -497 -1293 -481
rect -1235 -447 -1135 -400
rect -1235 -481 -1219 -447
rect -1151 -481 -1135 -447
rect -1235 -497 -1135 -481
rect -1077 -447 -977 -400
rect -1077 -481 -1061 -447
rect -993 -481 -977 -447
rect -1077 -497 -977 -481
rect -919 -447 -819 -400
rect -919 -481 -903 -447
rect -835 -481 -819 -447
rect -919 -497 -819 -481
rect -761 -447 -661 -400
rect -761 -481 -745 -447
rect -677 -481 -661 -447
rect -761 -497 -661 -481
rect -603 -447 -503 -400
rect -603 -481 -587 -447
rect -519 -481 -503 -447
rect -603 -497 -503 -481
rect -445 -447 -345 -400
rect -445 -481 -429 -447
rect -361 -481 -345 -447
rect -445 -497 -345 -481
rect -287 -447 -187 -400
rect -287 -481 -271 -447
rect -203 -481 -187 -447
rect -287 -497 -187 -481
rect -129 -447 -29 -400
rect -129 -481 -113 -447
rect -45 -481 -29 -447
rect -129 -497 -29 -481
rect 29 -447 129 -400
rect 29 -481 45 -447
rect 113 -481 129 -447
rect 29 -497 129 -481
rect 187 -447 287 -400
rect 187 -481 203 -447
rect 271 -481 287 -447
rect 187 -497 287 -481
rect 345 -447 445 -400
rect 345 -481 361 -447
rect 429 -481 445 -447
rect 345 -497 445 -481
rect 503 -447 603 -400
rect 503 -481 519 -447
rect 587 -481 603 -447
rect 503 -497 603 -481
rect 661 -447 761 -400
rect 661 -481 677 -447
rect 745 -481 761 -447
rect 661 -497 761 -481
rect 819 -447 919 -400
rect 819 -481 835 -447
rect 903 -481 919 -447
rect 819 -497 919 -481
rect 977 -447 1077 -400
rect 977 -481 993 -447
rect 1061 -481 1077 -447
rect 977 -497 1077 -481
rect 1135 -447 1235 -400
rect 1135 -481 1151 -447
rect 1219 -481 1235 -447
rect 1135 -497 1235 -481
rect 1293 -447 1393 -400
rect 1293 -481 1309 -447
rect 1377 -481 1393 -447
rect 1293 -497 1393 -481
rect 1451 -447 1551 -400
rect 1451 -481 1467 -447
rect 1535 -481 1551 -447
rect 1451 -497 1551 -481
rect 1609 -447 1709 -400
rect 1609 -481 1625 -447
rect 1693 -481 1709 -447
rect 1609 -497 1709 -481
rect 1767 -447 1867 -400
rect 1767 -481 1783 -447
rect 1851 -481 1867 -447
rect 1767 -497 1867 -481
rect 1925 -447 2025 -400
rect 1925 -481 1941 -447
rect 2009 -481 2025 -447
rect 1925 -497 2025 -481
rect 2083 -447 2183 -400
rect 2083 -481 2099 -447
rect 2167 -481 2183 -447
rect 2083 -497 2183 -481
rect 2241 -447 2341 -400
rect 2241 -481 2257 -447
rect 2325 -481 2341 -447
rect 2241 -497 2341 -481
rect 2399 -447 2499 -400
rect 2399 -481 2415 -447
rect 2483 -481 2499 -447
rect 2399 -497 2499 -481
rect 2557 -447 2657 -400
rect 2557 -481 2573 -447
rect 2641 -481 2657 -447
rect 2557 -497 2657 -481
rect 2715 -447 2815 -400
rect 2715 -481 2731 -447
rect 2799 -481 2815 -447
rect 2715 -497 2815 -481
rect 2873 -447 2973 -400
rect 2873 -481 2889 -447
rect 2957 -481 2973 -447
rect 2873 -497 2973 -481
rect 3031 -447 3131 -400
rect 3031 -481 3047 -447
rect 3115 -481 3131 -447
rect 3031 -497 3131 -481
rect 3189 -447 3289 -400
rect 3189 -481 3205 -447
rect 3273 -481 3289 -447
rect 3189 -497 3289 -481
rect 3347 -447 3447 -400
rect 3347 -481 3363 -447
rect 3431 -481 3447 -447
rect 3347 -497 3447 -481
rect 3505 -447 3605 -400
rect 3505 -481 3521 -447
rect 3589 -481 3605 -447
rect 3505 -497 3605 -481
rect 3663 -447 3763 -400
rect 3663 -481 3679 -447
rect 3747 -481 3763 -447
rect 3663 -497 3763 -481
rect 3821 -447 3921 -400
rect 3821 -481 3837 -447
rect 3905 -481 3921 -447
rect 3821 -497 3921 -481
rect 3979 -447 4079 -400
rect 3979 -481 3995 -447
rect 4063 -481 4079 -447
rect 3979 -497 4079 -481
rect 4137 -447 4237 -400
rect 4137 -481 4153 -447
rect 4221 -481 4237 -447
rect 4137 -497 4237 -481
rect 4295 -447 4395 -400
rect 4295 -481 4311 -447
rect 4379 -481 4395 -447
rect 4295 -497 4395 -481
rect 4453 -447 4553 -400
rect 4453 -481 4469 -447
rect 4537 -481 4553 -447
rect 4453 -497 4553 -481
rect 4611 -447 4711 -400
rect 4611 -481 4627 -447
rect 4695 -481 4711 -447
rect 4611 -497 4711 -481
rect 4769 -447 4869 -400
rect 4769 -481 4785 -447
rect 4853 -481 4869 -447
rect 4769 -497 4869 -481
rect 4927 -447 5027 -400
rect 4927 -481 4943 -447
rect 5011 -481 5027 -447
rect 4927 -497 5027 -481
rect 5085 -447 5185 -400
rect 5085 -481 5101 -447
rect 5169 -481 5185 -447
rect 5085 -497 5185 -481
rect 5243 -447 5343 -400
rect 5243 -481 5259 -447
rect 5327 -481 5343 -447
rect 5243 -497 5343 -481
rect 5401 -447 5501 -400
rect 5401 -481 5417 -447
rect 5485 -481 5501 -447
rect 5401 -497 5501 -481
rect 5559 -447 5659 -400
rect 5559 -481 5575 -447
rect 5643 -481 5659 -447
rect 5559 -497 5659 -481
rect 5717 -447 5817 -400
rect 5717 -481 5733 -447
rect 5801 -481 5817 -447
rect 5717 -497 5817 -481
rect 5875 -447 5975 -400
rect 5875 -481 5891 -447
rect 5959 -481 5975 -447
rect 5875 -497 5975 -481
rect 6033 -447 6133 -400
rect 6033 -481 6049 -447
rect 6117 -481 6133 -447
rect 6033 -497 6133 -481
rect 6191 -447 6291 -400
rect 6191 -481 6207 -447
rect 6275 -481 6291 -447
rect 6191 -497 6291 -481
<< polycont >>
rect -6275 447 -6207 481
rect -6117 447 -6049 481
rect -5959 447 -5891 481
rect -5801 447 -5733 481
rect -5643 447 -5575 481
rect -5485 447 -5417 481
rect -5327 447 -5259 481
rect -5169 447 -5101 481
rect -5011 447 -4943 481
rect -4853 447 -4785 481
rect -4695 447 -4627 481
rect -4537 447 -4469 481
rect -4379 447 -4311 481
rect -4221 447 -4153 481
rect -4063 447 -3995 481
rect -3905 447 -3837 481
rect -3747 447 -3679 481
rect -3589 447 -3521 481
rect -3431 447 -3363 481
rect -3273 447 -3205 481
rect -3115 447 -3047 481
rect -2957 447 -2889 481
rect -2799 447 -2731 481
rect -2641 447 -2573 481
rect -2483 447 -2415 481
rect -2325 447 -2257 481
rect -2167 447 -2099 481
rect -2009 447 -1941 481
rect -1851 447 -1783 481
rect -1693 447 -1625 481
rect -1535 447 -1467 481
rect -1377 447 -1309 481
rect -1219 447 -1151 481
rect -1061 447 -993 481
rect -903 447 -835 481
rect -745 447 -677 481
rect -587 447 -519 481
rect -429 447 -361 481
rect -271 447 -203 481
rect -113 447 -45 481
rect 45 447 113 481
rect 203 447 271 481
rect 361 447 429 481
rect 519 447 587 481
rect 677 447 745 481
rect 835 447 903 481
rect 993 447 1061 481
rect 1151 447 1219 481
rect 1309 447 1377 481
rect 1467 447 1535 481
rect 1625 447 1693 481
rect 1783 447 1851 481
rect 1941 447 2009 481
rect 2099 447 2167 481
rect 2257 447 2325 481
rect 2415 447 2483 481
rect 2573 447 2641 481
rect 2731 447 2799 481
rect 2889 447 2957 481
rect 3047 447 3115 481
rect 3205 447 3273 481
rect 3363 447 3431 481
rect 3521 447 3589 481
rect 3679 447 3747 481
rect 3837 447 3905 481
rect 3995 447 4063 481
rect 4153 447 4221 481
rect 4311 447 4379 481
rect 4469 447 4537 481
rect 4627 447 4695 481
rect 4785 447 4853 481
rect 4943 447 5011 481
rect 5101 447 5169 481
rect 5259 447 5327 481
rect 5417 447 5485 481
rect 5575 447 5643 481
rect 5733 447 5801 481
rect 5891 447 5959 481
rect 6049 447 6117 481
rect 6207 447 6275 481
rect -6275 -481 -6207 -447
rect -6117 -481 -6049 -447
rect -5959 -481 -5891 -447
rect -5801 -481 -5733 -447
rect -5643 -481 -5575 -447
rect -5485 -481 -5417 -447
rect -5327 -481 -5259 -447
rect -5169 -481 -5101 -447
rect -5011 -481 -4943 -447
rect -4853 -481 -4785 -447
rect -4695 -481 -4627 -447
rect -4537 -481 -4469 -447
rect -4379 -481 -4311 -447
rect -4221 -481 -4153 -447
rect -4063 -481 -3995 -447
rect -3905 -481 -3837 -447
rect -3747 -481 -3679 -447
rect -3589 -481 -3521 -447
rect -3431 -481 -3363 -447
rect -3273 -481 -3205 -447
rect -3115 -481 -3047 -447
rect -2957 -481 -2889 -447
rect -2799 -481 -2731 -447
rect -2641 -481 -2573 -447
rect -2483 -481 -2415 -447
rect -2325 -481 -2257 -447
rect -2167 -481 -2099 -447
rect -2009 -481 -1941 -447
rect -1851 -481 -1783 -447
rect -1693 -481 -1625 -447
rect -1535 -481 -1467 -447
rect -1377 -481 -1309 -447
rect -1219 -481 -1151 -447
rect -1061 -481 -993 -447
rect -903 -481 -835 -447
rect -745 -481 -677 -447
rect -587 -481 -519 -447
rect -429 -481 -361 -447
rect -271 -481 -203 -447
rect -113 -481 -45 -447
rect 45 -481 113 -447
rect 203 -481 271 -447
rect 361 -481 429 -447
rect 519 -481 587 -447
rect 677 -481 745 -447
rect 835 -481 903 -447
rect 993 -481 1061 -447
rect 1151 -481 1219 -447
rect 1309 -481 1377 -447
rect 1467 -481 1535 -447
rect 1625 -481 1693 -447
rect 1783 -481 1851 -447
rect 1941 -481 2009 -447
rect 2099 -481 2167 -447
rect 2257 -481 2325 -447
rect 2415 -481 2483 -447
rect 2573 -481 2641 -447
rect 2731 -481 2799 -447
rect 2889 -481 2957 -447
rect 3047 -481 3115 -447
rect 3205 -481 3273 -447
rect 3363 -481 3431 -447
rect 3521 -481 3589 -447
rect 3679 -481 3747 -447
rect 3837 -481 3905 -447
rect 3995 -481 4063 -447
rect 4153 -481 4221 -447
rect 4311 -481 4379 -447
rect 4469 -481 4537 -447
rect 4627 -481 4695 -447
rect 4785 -481 4853 -447
rect 4943 -481 5011 -447
rect 5101 -481 5169 -447
rect 5259 -481 5327 -447
rect 5417 -481 5485 -447
rect 5575 -481 5643 -447
rect 5733 -481 5801 -447
rect 5891 -481 5959 -447
rect 6049 -481 6117 -447
rect 6207 -481 6275 -447
<< locali >>
rect -6471 585 -6375 619
rect 6375 585 6471 619
rect -6471 523 -6437 585
rect 6437 523 6471 585
rect -6291 447 -6275 481
rect -6207 447 -6191 481
rect -6133 447 -6117 481
rect -6049 447 -6033 481
rect -5975 447 -5959 481
rect -5891 447 -5875 481
rect -5817 447 -5801 481
rect -5733 447 -5717 481
rect -5659 447 -5643 481
rect -5575 447 -5559 481
rect -5501 447 -5485 481
rect -5417 447 -5401 481
rect -5343 447 -5327 481
rect -5259 447 -5243 481
rect -5185 447 -5169 481
rect -5101 447 -5085 481
rect -5027 447 -5011 481
rect -4943 447 -4927 481
rect -4869 447 -4853 481
rect -4785 447 -4769 481
rect -4711 447 -4695 481
rect -4627 447 -4611 481
rect -4553 447 -4537 481
rect -4469 447 -4453 481
rect -4395 447 -4379 481
rect -4311 447 -4295 481
rect -4237 447 -4221 481
rect -4153 447 -4137 481
rect -4079 447 -4063 481
rect -3995 447 -3979 481
rect -3921 447 -3905 481
rect -3837 447 -3821 481
rect -3763 447 -3747 481
rect -3679 447 -3663 481
rect -3605 447 -3589 481
rect -3521 447 -3505 481
rect -3447 447 -3431 481
rect -3363 447 -3347 481
rect -3289 447 -3273 481
rect -3205 447 -3189 481
rect -3131 447 -3115 481
rect -3047 447 -3031 481
rect -2973 447 -2957 481
rect -2889 447 -2873 481
rect -2815 447 -2799 481
rect -2731 447 -2715 481
rect -2657 447 -2641 481
rect -2573 447 -2557 481
rect -2499 447 -2483 481
rect -2415 447 -2399 481
rect -2341 447 -2325 481
rect -2257 447 -2241 481
rect -2183 447 -2167 481
rect -2099 447 -2083 481
rect -2025 447 -2009 481
rect -1941 447 -1925 481
rect -1867 447 -1851 481
rect -1783 447 -1767 481
rect -1709 447 -1693 481
rect -1625 447 -1609 481
rect -1551 447 -1535 481
rect -1467 447 -1451 481
rect -1393 447 -1377 481
rect -1309 447 -1293 481
rect -1235 447 -1219 481
rect -1151 447 -1135 481
rect -1077 447 -1061 481
rect -993 447 -977 481
rect -919 447 -903 481
rect -835 447 -819 481
rect -761 447 -745 481
rect -677 447 -661 481
rect -603 447 -587 481
rect -519 447 -503 481
rect -445 447 -429 481
rect -361 447 -345 481
rect -287 447 -271 481
rect -203 447 -187 481
rect -129 447 -113 481
rect -45 447 -29 481
rect 29 447 45 481
rect 113 447 129 481
rect 187 447 203 481
rect 271 447 287 481
rect 345 447 361 481
rect 429 447 445 481
rect 503 447 519 481
rect 587 447 603 481
rect 661 447 677 481
rect 745 447 761 481
rect 819 447 835 481
rect 903 447 919 481
rect 977 447 993 481
rect 1061 447 1077 481
rect 1135 447 1151 481
rect 1219 447 1235 481
rect 1293 447 1309 481
rect 1377 447 1393 481
rect 1451 447 1467 481
rect 1535 447 1551 481
rect 1609 447 1625 481
rect 1693 447 1709 481
rect 1767 447 1783 481
rect 1851 447 1867 481
rect 1925 447 1941 481
rect 2009 447 2025 481
rect 2083 447 2099 481
rect 2167 447 2183 481
rect 2241 447 2257 481
rect 2325 447 2341 481
rect 2399 447 2415 481
rect 2483 447 2499 481
rect 2557 447 2573 481
rect 2641 447 2657 481
rect 2715 447 2731 481
rect 2799 447 2815 481
rect 2873 447 2889 481
rect 2957 447 2973 481
rect 3031 447 3047 481
rect 3115 447 3131 481
rect 3189 447 3205 481
rect 3273 447 3289 481
rect 3347 447 3363 481
rect 3431 447 3447 481
rect 3505 447 3521 481
rect 3589 447 3605 481
rect 3663 447 3679 481
rect 3747 447 3763 481
rect 3821 447 3837 481
rect 3905 447 3921 481
rect 3979 447 3995 481
rect 4063 447 4079 481
rect 4137 447 4153 481
rect 4221 447 4237 481
rect 4295 447 4311 481
rect 4379 447 4395 481
rect 4453 447 4469 481
rect 4537 447 4553 481
rect 4611 447 4627 481
rect 4695 447 4711 481
rect 4769 447 4785 481
rect 4853 447 4869 481
rect 4927 447 4943 481
rect 5011 447 5027 481
rect 5085 447 5101 481
rect 5169 447 5185 481
rect 5243 447 5259 481
rect 5327 447 5343 481
rect 5401 447 5417 481
rect 5485 447 5501 481
rect 5559 447 5575 481
rect 5643 447 5659 481
rect 5717 447 5733 481
rect 5801 447 5817 481
rect 5875 447 5891 481
rect 5959 447 5975 481
rect 6033 447 6049 481
rect 6117 447 6133 481
rect 6191 447 6207 481
rect 6275 447 6291 481
rect -6337 388 -6303 404
rect -6337 -404 -6303 -388
rect -6179 388 -6145 404
rect -6179 -404 -6145 -388
rect -6021 388 -5987 404
rect -6021 -404 -5987 -388
rect -5863 388 -5829 404
rect -5863 -404 -5829 -388
rect -5705 388 -5671 404
rect -5705 -404 -5671 -388
rect -5547 388 -5513 404
rect -5547 -404 -5513 -388
rect -5389 388 -5355 404
rect -5389 -404 -5355 -388
rect -5231 388 -5197 404
rect -5231 -404 -5197 -388
rect -5073 388 -5039 404
rect -5073 -404 -5039 -388
rect -4915 388 -4881 404
rect -4915 -404 -4881 -388
rect -4757 388 -4723 404
rect -4757 -404 -4723 -388
rect -4599 388 -4565 404
rect -4599 -404 -4565 -388
rect -4441 388 -4407 404
rect -4441 -404 -4407 -388
rect -4283 388 -4249 404
rect -4283 -404 -4249 -388
rect -4125 388 -4091 404
rect -4125 -404 -4091 -388
rect -3967 388 -3933 404
rect -3967 -404 -3933 -388
rect -3809 388 -3775 404
rect -3809 -404 -3775 -388
rect -3651 388 -3617 404
rect -3651 -404 -3617 -388
rect -3493 388 -3459 404
rect -3493 -404 -3459 -388
rect -3335 388 -3301 404
rect -3335 -404 -3301 -388
rect -3177 388 -3143 404
rect -3177 -404 -3143 -388
rect -3019 388 -2985 404
rect -3019 -404 -2985 -388
rect -2861 388 -2827 404
rect -2861 -404 -2827 -388
rect -2703 388 -2669 404
rect -2703 -404 -2669 -388
rect -2545 388 -2511 404
rect -2545 -404 -2511 -388
rect -2387 388 -2353 404
rect -2387 -404 -2353 -388
rect -2229 388 -2195 404
rect -2229 -404 -2195 -388
rect -2071 388 -2037 404
rect -2071 -404 -2037 -388
rect -1913 388 -1879 404
rect -1913 -404 -1879 -388
rect -1755 388 -1721 404
rect -1755 -404 -1721 -388
rect -1597 388 -1563 404
rect -1597 -404 -1563 -388
rect -1439 388 -1405 404
rect -1439 -404 -1405 -388
rect -1281 388 -1247 404
rect -1281 -404 -1247 -388
rect -1123 388 -1089 404
rect -1123 -404 -1089 -388
rect -965 388 -931 404
rect -965 -404 -931 -388
rect -807 388 -773 404
rect -807 -404 -773 -388
rect -649 388 -615 404
rect -649 -404 -615 -388
rect -491 388 -457 404
rect -491 -404 -457 -388
rect -333 388 -299 404
rect -333 -404 -299 -388
rect -175 388 -141 404
rect -175 -404 -141 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 141 388 175 404
rect 141 -404 175 -388
rect 299 388 333 404
rect 299 -404 333 -388
rect 457 388 491 404
rect 457 -404 491 -388
rect 615 388 649 404
rect 615 -404 649 -388
rect 773 388 807 404
rect 773 -404 807 -388
rect 931 388 965 404
rect 931 -404 965 -388
rect 1089 388 1123 404
rect 1089 -404 1123 -388
rect 1247 388 1281 404
rect 1247 -404 1281 -388
rect 1405 388 1439 404
rect 1405 -404 1439 -388
rect 1563 388 1597 404
rect 1563 -404 1597 -388
rect 1721 388 1755 404
rect 1721 -404 1755 -388
rect 1879 388 1913 404
rect 1879 -404 1913 -388
rect 2037 388 2071 404
rect 2037 -404 2071 -388
rect 2195 388 2229 404
rect 2195 -404 2229 -388
rect 2353 388 2387 404
rect 2353 -404 2387 -388
rect 2511 388 2545 404
rect 2511 -404 2545 -388
rect 2669 388 2703 404
rect 2669 -404 2703 -388
rect 2827 388 2861 404
rect 2827 -404 2861 -388
rect 2985 388 3019 404
rect 2985 -404 3019 -388
rect 3143 388 3177 404
rect 3143 -404 3177 -388
rect 3301 388 3335 404
rect 3301 -404 3335 -388
rect 3459 388 3493 404
rect 3459 -404 3493 -388
rect 3617 388 3651 404
rect 3617 -404 3651 -388
rect 3775 388 3809 404
rect 3775 -404 3809 -388
rect 3933 388 3967 404
rect 3933 -404 3967 -388
rect 4091 388 4125 404
rect 4091 -404 4125 -388
rect 4249 388 4283 404
rect 4249 -404 4283 -388
rect 4407 388 4441 404
rect 4407 -404 4441 -388
rect 4565 388 4599 404
rect 4565 -404 4599 -388
rect 4723 388 4757 404
rect 4723 -404 4757 -388
rect 4881 388 4915 404
rect 4881 -404 4915 -388
rect 5039 388 5073 404
rect 5039 -404 5073 -388
rect 5197 388 5231 404
rect 5197 -404 5231 -388
rect 5355 388 5389 404
rect 5355 -404 5389 -388
rect 5513 388 5547 404
rect 5513 -404 5547 -388
rect 5671 388 5705 404
rect 5671 -404 5705 -388
rect 5829 388 5863 404
rect 5829 -404 5863 -388
rect 5987 388 6021 404
rect 5987 -404 6021 -388
rect 6145 388 6179 404
rect 6145 -404 6179 -388
rect 6303 388 6337 404
rect 6303 -404 6337 -388
rect -6291 -481 -6275 -447
rect -6207 -481 -6191 -447
rect -6133 -481 -6117 -447
rect -6049 -481 -6033 -447
rect -5975 -481 -5959 -447
rect -5891 -481 -5875 -447
rect -5817 -481 -5801 -447
rect -5733 -481 -5717 -447
rect -5659 -481 -5643 -447
rect -5575 -481 -5559 -447
rect -5501 -481 -5485 -447
rect -5417 -481 -5401 -447
rect -5343 -481 -5327 -447
rect -5259 -481 -5243 -447
rect -5185 -481 -5169 -447
rect -5101 -481 -5085 -447
rect -5027 -481 -5011 -447
rect -4943 -481 -4927 -447
rect -4869 -481 -4853 -447
rect -4785 -481 -4769 -447
rect -4711 -481 -4695 -447
rect -4627 -481 -4611 -447
rect -4553 -481 -4537 -447
rect -4469 -481 -4453 -447
rect -4395 -481 -4379 -447
rect -4311 -481 -4295 -447
rect -4237 -481 -4221 -447
rect -4153 -481 -4137 -447
rect -4079 -481 -4063 -447
rect -3995 -481 -3979 -447
rect -3921 -481 -3905 -447
rect -3837 -481 -3821 -447
rect -3763 -481 -3747 -447
rect -3679 -481 -3663 -447
rect -3605 -481 -3589 -447
rect -3521 -481 -3505 -447
rect -3447 -481 -3431 -447
rect -3363 -481 -3347 -447
rect -3289 -481 -3273 -447
rect -3205 -481 -3189 -447
rect -3131 -481 -3115 -447
rect -3047 -481 -3031 -447
rect -2973 -481 -2957 -447
rect -2889 -481 -2873 -447
rect -2815 -481 -2799 -447
rect -2731 -481 -2715 -447
rect -2657 -481 -2641 -447
rect -2573 -481 -2557 -447
rect -2499 -481 -2483 -447
rect -2415 -481 -2399 -447
rect -2341 -481 -2325 -447
rect -2257 -481 -2241 -447
rect -2183 -481 -2167 -447
rect -2099 -481 -2083 -447
rect -2025 -481 -2009 -447
rect -1941 -481 -1925 -447
rect -1867 -481 -1851 -447
rect -1783 -481 -1767 -447
rect -1709 -481 -1693 -447
rect -1625 -481 -1609 -447
rect -1551 -481 -1535 -447
rect -1467 -481 -1451 -447
rect -1393 -481 -1377 -447
rect -1309 -481 -1293 -447
rect -1235 -481 -1219 -447
rect -1151 -481 -1135 -447
rect -1077 -481 -1061 -447
rect -993 -481 -977 -447
rect -919 -481 -903 -447
rect -835 -481 -819 -447
rect -761 -481 -745 -447
rect -677 -481 -661 -447
rect -603 -481 -587 -447
rect -519 -481 -503 -447
rect -445 -481 -429 -447
rect -361 -481 -345 -447
rect -287 -481 -271 -447
rect -203 -481 -187 -447
rect -129 -481 -113 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 113 -481 129 -447
rect 187 -481 203 -447
rect 271 -481 287 -447
rect 345 -481 361 -447
rect 429 -481 445 -447
rect 503 -481 519 -447
rect 587 -481 603 -447
rect 661 -481 677 -447
rect 745 -481 761 -447
rect 819 -481 835 -447
rect 903 -481 919 -447
rect 977 -481 993 -447
rect 1061 -481 1077 -447
rect 1135 -481 1151 -447
rect 1219 -481 1235 -447
rect 1293 -481 1309 -447
rect 1377 -481 1393 -447
rect 1451 -481 1467 -447
rect 1535 -481 1551 -447
rect 1609 -481 1625 -447
rect 1693 -481 1709 -447
rect 1767 -481 1783 -447
rect 1851 -481 1867 -447
rect 1925 -481 1941 -447
rect 2009 -481 2025 -447
rect 2083 -481 2099 -447
rect 2167 -481 2183 -447
rect 2241 -481 2257 -447
rect 2325 -481 2341 -447
rect 2399 -481 2415 -447
rect 2483 -481 2499 -447
rect 2557 -481 2573 -447
rect 2641 -481 2657 -447
rect 2715 -481 2731 -447
rect 2799 -481 2815 -447
rect 2873 -481 2889 -447
rect 2957 -481 2973 -447
rect 3031 -481 3047 -447
rect 3115 -481 3131 -447
rect 3189 -481 3205 -447
rect 3273 -481 3289 -447
rect 3347 -481 3363 -447
rect 3431 -481 3447 -447
rect 3505 -481 3521 -447
rect 3589 -481 3605 -447
rect 3663 -481 3679 -447
rect 3747 -481 3763 -447
rect 3821 -481 3837 -447
rect 3905 -481 3921 -447
rect 3979 -481 3995 -447
rect 4063 -481 4079 -447
rect 4137 -481 4153 -447
rect 4221 -481 4237 -447
rect 4295 -481 4311 -447
rect 4379 -481 4395 -447
rect 4453 -481 4469 -447
rect 4537 -481 4553 -447
rect 4611 -481 4627 -447
rect 4695 -481 4711 -447
rect 4769 -481 4785 -447
rect 4853 -481 4869 -447
rect 4927 -481 4943 -447
rect 5011 -481 5027 -447
rect 5085 -481 5101 -447
rect 5169 -481 5185 -447
rect 5243 -481 5259 -447
rect 5327 -481 5343 -447
rect 5401 -481 5417 -447
rect 5485 -481 5501 -447
rect 5559 -481 5575 -447
rect 5643 -481 5659 -447
rect 5717 -481 5733 -447
rect 5801 -481 5817 -447
rect 5875 -481 5891 -447
rect 5959 -481 5975 -447
rect 6033 -481 6049 -447
rect 6117 -481 6133 -447
rect 6191 -481 6207 -447
rect 6275 -481 6291 -447
rect -6471 -585 -6437 -523
rect 6437 -585 6471 -523
rect -6471 -619 -6375 -585
rect 6375 -619 6471 -585
<< viali >>
rect -6275 447 -6207 481
rect -6117 447 -6049 481
rect -5959 447 -5891 481
rect -5801 447 -5733 481
rect -5643 447 -5575 481
rect -5485 447 -5417 481
rect -5327 447 -5259 481
rect -5169 447 -5101 481
rect -5011 447 -4943 481
rect -4853 447 -4785 481
rect -4695 447 -4627 481
rect -4537 447 -4469 481
rect -4379 447 -4311 481
rect -4221 447 -4153 481
rect -4063 447 -3995 481
rect -3905 447 -3837 481
rect -3747 447 -3679 481
rect -3589 447 -3521 481
rect -3431 447 -3363 481
rect -3273 447 -3205 481
rect -3115 447 -3047 481
rect -2957 447 -2889 481
rect -2799 447 -2731 481
rect -2641 447 -2573 481
rect -2483 447 -2415 481
rect -2325 447 -2257 481
rect -2167 447 -2099 481
rect -2009 447 -1941 481
rect -1851 447 -1783 481
rect -1693 447 -1625 481
rect -1535 447 -1467 481
rect -1377 447 -1309 481
rect -1219 447 -1151 481
rect -1061 447 -993 481
rect -903 447 -835 481
rect -745 447 -677 481
rect -587 447 -519 481
rect -429 447 -361 481
rect -271 447 -203 481
rect -113 447 -45 481
rect 45 447 113 481
rect 203 447 271 481
rect 361 447 429 481
rect 519 447 587 481
rect 677 447 745 481
rect 835 447 903 481
rect 993 447 1061 481
rect 1151 447 1219 481
rect 1309 447 1377 481
rect 1467 447 1535 481
rect 1625 447 1693 481
rect 1783 447 1851 481
rect 1941 447 2009 481
rect 2099 447 2167 481
rect 2257 447 2325 481
rect 2415 447 2483 481
rect 2573 447 2641 481
rect 2731 447 2799 481
rect 2889 447 2957 481
rect 3047 447 3115 481
rect 3205 447 3273 481
rect 3363 447 3431 481
rect 3521 447 3589 481
rect 3679 447 3747 481
rect 3837 447 3905 481
rect 3995 447 4063 481
rect 4153 447 4221 481
rect 4311 447 4379 481
rect 4469 447 4537 481
rect 4627 447 4695 481
rect 4785 447 4853 481
rect 4943 447 5011 481
rect 5101 447 5169 481
rect 5259 447 5327 481
rect 5417 447 5485 481
rect 5575 447 5643 481
rect 5733 447 5801 481
rect 5891 447 5959 481
rect 6049 447 6117 481
rect 6207 447 6275 481
rect -6337 -388 -6303 388
rect -6179 -388 -6145 388
rect -6021 -388 -5987 388
rect -5863 -388 -5829 388
rect -5705 -388 -5671 388
rect -5547 -388 -5513 388
rect -5389 -388 -5355 388
rect -5231 -388 -5197 388
rect -5073 -388 -5039 388
rect -4915 -388 -4881 388
rect -4757 -388 -4723 388
rect -4599 -388 -4565 388
rect -4441 -388 -4407 388
rect -4283 -388 -4249 388
rect -4125 -388 -4091 388
rect -3967 -388 -3933 388
rect -3809 -388 -3775 388
rect -3651 -388 -3617 388
rect -3493 -388 -3459 388
rect -3335 -388 -3301 388
rect -3177 -388 -3143 388
rect -3019 -388 -2985 388
rect -2861 -388 -2827 388
rect -2703 -388 -2669 388
rect -2545 -388 -2511 388
rect -2387 -388 -2353 388
rect -2229 -388 -2195 388
rect -2071 -388 -2037 388
rect -1913 -388 -1879 388
rect -1755 -388 -1721 388
rect -1597 -388 -1563 388
rect -1439 -388 -1405 388
rect -1281 -388 -1247 388
rect -1123 -388 -1089 388
rect -965 -388 -931 388
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
rect 931 -388 965 388
rect 1089 -388 1123 388
rect 1247 -388 1281 388
rect 1405 -388 1439 388
rect 1563 -388 1597 388
rect 1721 -388 1755 388
rect 1879 -388 1913 388
rect 2037 -388 2071 388
rect 2195 -388 2229 388
rect 2353 -388 2387 388
rect 2511 -388 2545 388
rect 2669 -388 2703 388
rect 2827 -388 2861 388
rect 2985 -388 3019 388
rect 3143 -388 3177 388
rect 3301 -388 3335 388
rect 3459 -388 3493 388
rect 3617 -388 3651 388
rect 3775 -388 3809 388
rect 3933 -388 3967 388
rect 4091 -388 4125 388
rect 4249 -388 4283 388
rect 4407 -388 4441 388
rect 4565 -388 4599 388
rect 4723 -388 4757 388
rect 4881 -388 4915 388
rect 5039 -388 5073 388
rect 5197 -388 5231 388
rect 5355 -388 5389 388
rect 5513 -388 5547 388
rect 5671 -388 5705 388
rect 5829 -388 5863 388
rect 5987 -388 6021 388
rect 6145 -388 6179 388
rect 6303 -388 6337 388
rect -6275 -481 -6207 -447
rect -6117 -481 -6049 -447
rect -5959 -481 -5891 -447
rect -5801 -481 -5733 -447
rect -5643 -481 -5575 -447
rect -5485 -481 -5417 -447
rect -5327 -481 -5259 -447
rect -5169 -481 -5101 -447
rect -5011 -481 -4943 -447
rect -4853 -481 -4785 -447
rect -4695 -481 -4627 -447
rect -4537 -481 -4469 -447
rect -4379 -481 -4311 -447
rect -4221 -481 -4153 -447
rect -4063 -481 -3995 -447
rect -3905 -481 -3837 -447
rect -3747 -481 -3679 -447
rect -3589 -481 -3521 -447
rect -3431 -481 -3363 -447
rect -3273 -481 -3205 -447
rect -3115 -481 -3047 -447
rect -2957 -481 -2889 -447
rect -2799 -481 -2731 -447
rect -2641 -481 -2573 -447
rect -2483 -481 -2415 -447
rect -2325 -481 -2257 -447
rect -2167 -481 -2099 -447
rect -2009 -481 -1941 -447
rect -1851 -481 -1783 -447
rect -1693 -481 -1625 -447
rect -1535 -481 -1467 -447
rect -1377 -481 -1309 -447
rect -1219 -481 -1151 -447
rect -1061 -481 -993 -447
rect -903 -481 -835 -447
rect -745 -481 -677 -447
rect -587 -481 -519 -447
rect -429 -481 -361 -447
rect -271 -481 -203 -447
rect -113 -481 -45 -447
rect 45 -481 113 -447
rect 203 -481 271 -447
rect 361 -481 429 -447
rect 519 -481 587 -447
rect 677 -481 745 -447
rect 835 -481 903 -447
rect 993 -481 1061 -447
rect 1151 -481 1219 -447
rect 1309 -481 1377 -447
rect 1467 -481 1535 -447
rect 1625 -481 1693 -447
rect 1783 -481 1851 -447
rect 1941 -481 2009 -447
rect 2099 -481 2167 -447
rect 2257 -481 2325 -447
rect 2415 -481 2483 -447
rect 2573 -481 2641 -447
rect 2731 -481 2799 -447
rect 2889 -481 2957 -447
rect 3047 -481 3115 -447
rect 3205 -481 3273 -447
rect 3363 -481 3431 -447
rect 3521 -481 3589 -447
rect 3679 -481 3747 -447
rect 3837 -481 3905 -447
rect 3995 -481 4063 -447
rect 4153 -481 4221 -447
rect 4311 -481 4379 -447
rect 4469 -481 4537 -447
rect 4627 -481 4695 -447
rect 4785 -481 4853 -447
rect 4943 -481 5011 -447
rect 5101 -481 5169 -447
rect 5259 -481 5327 -447
rect 5417 -481 5485 -447
rect 5575 -481 5643 -447
rect 5733 -481 5801 -447
rect 5891 -481 5959 -447
rect 6049 -481 6117 -447
rect 6207 -481 6275 -447
<< metal1 >>
rect -6287 481 -6195 487
rect -6287 447 -6275 481
rect -6207 447 -6195 481
rect -6287 441 -6195 447
rect -6129 481 -6037 487
rect -6129 447 -6117 481
rect -6049 447 -6037 481
rect -6129 441 -6037 447
rect -5971 481 -5879 487
rect -5971 447 -5959 481
rect -5891 447 -5879 481
rect -5971 441 -5879 447
rect -5813 481 -5721 487
rect -5813 447 -5801 481
rect -5733 447 -5721 481
rect -5813 441 -5721 447
rect -5655 481 -5563 487
rect -5655 447 -5643 481
rect -5575 447 -5563 481
rect -5655 441 -5563 447
rect -5497 481 -5405 487
rect -5497 447 -5485 481
rect -5417 447 -5405 481
rect -5497 441 -5405 447
rect -5339 481 -5247 487
rect -5339 447 -5327 481
rect -5259 447 -5247 481
rect -5339 441 -5247 447
rect -5181 481 -5089 487
rect -5181 447 -5169 481
rect -5101 447 -5089 481
rect -5181 441 -5089 447
rect -5023 481 -4931 487
rect -5023 447 -5011 481
rect -4943 447 -4931 481
rect -5023 441 -4931 447
rect -4865 481 -4773 487
rect -4865 447 -4853 481
rect -4785 447 -4773 481
rect -4865 441 -4773 447
rect -4707 481 -4615 487
rect -4707 447 -4695 481
rect -4627 447 -4615 481
rect -4707 441 -4615 447
rect -4549 481 -4457 487
rect -4549 447 -4537 481
rect -4469 447 -4457 481
rect -4549 441 -4457 447
rect -4391 481 -4299 487
rect -4391 447 -4379 481
rect -4311 447 -4299 481
rect -4391 441 -4299 447
rect -4233 481 -4141 487
rect -4233 447 -4221 481
rect -4153 447 -4141 481
rect -4233 441 -4141 447
rect -4075 481 -3983 487
rect -4075 447 -4063 481
rect -3995 447 -3983 481
rect -4075 441 -3983 447
rect -3917 481 -3825 487
rect -3917 447 -3905 481
rect -3837 447 -3825 481
rect -3917 441 -3825 447
rect -3759 481 -3667 487
rect -3759 447 -3747 481
rect -3679 447 -3667 481
rect -3759 441 -3667 447
rect -3601 481 -3509 487
rect -3601 447 -3589 481
rect -3521 447 -3509 481
rect -3601 441 -3509 447
rect -3443 481 -3351 487
rect -3443 447 -3431 481
rect -3363 447 -3351 481
rect -3443 441 -3351 447
rect -3285 481 -3193 487
rect -3285 447 -3273 481
rect -3205 447 -3193 481
rect -3285 441 -3193 447
rect -3127 481 -3035 487
rect -3127 447 -3115 481
rect -3047 447 -3035 481
rect -3127 441 -3035 447
rect -2969 481 -2877 487
rect -2969 447 -2957 481
rect -2889 447 -2877 481
rect -2969 441 -2877 447
rect -2811 481 -2719 487
rect -2811 447 -2799 481
rect -2731 447 -2719 481
rect -2811 441 -2719 447
rect -2653 481 -2561 487
rect -2653 447 -2641 481
rect -2573 447 -2561 481
rect -2653 441 -2561 447
rect -2495 481 -2403 487
rect -2495 447 -2483 481
rect -2415 447 -2403 481
rect -2495 441 -2403 447
rect -2337 481 -2245 487
rect -2337 447 -2325 481
rect -2257 447 -2245 481
rect -2337 441 -2245 447
rect -2179 481 -2087 487
rect -2179 447 -2167 481
rect -2099 447 -2087 481
rect -2179 441 -2087 447
rect -2021 481 -1929 487
rect -2021 447 -2009 481
rect -1941 447 -1929 481
rect -2021 441 -1929 447
rect -1863 481 -1771 487
rect -1863 447 -1851 481
rect -1783 447 -1771 481
rect -1863 441 -1771 447
rect -1705 481 -1613 487
rect -1705 447 -1693 481
rect -1625 447 -1613 481
rect -1705 441 -1613 447
rect -1547 481 -1455 487
rect -1547 447 -1535 481
rect -1467 447 -1455 481
rect -1547 441 -1455 447
rect -1389 481 -1297 487
rect -1389 447 -1377 481
rect -1309 447 -1297 481
rect -1389 441 -1297 447
rect -1231 481 -1139 487
rect -1231 447 -1219 481
rect -1151 447 -1139 481
rect -1231 441 -1139 447
rect -1073 481 -981 487
rect -1073 447 -1061 481
rect -993 447 -981 481
rect -1073 441 -981 447
rect -915 481 -823 487
rect -915 447 -903 481
rect -835 447 -823 481
rect -915 441 -823 447
rect -757 481 -665 487
rect -757 447 -745 481
rect -677 447 -665 481
rect -757 441 -665 447
rect -599 481 -507 487
rect -599 447 -587 481
rect -519 447 -507 481
rect -599 441 -507 447
rect -441 481 -349 487
rect -441 447 -429 481
rect -361 447 -349 481
rect -441 441 -349 447
rect -283 481 -191 487
rect -283 447 -271 481
rect -203 447 -191 481
rect -283 441 -191 447
rect -125 481 -33 487
rect -125 447 -113 481
rect -45 447 -33 481
rect -125 441 -33 447
rect 33 481 125 487
rect 33 447 45 481
rect 113 447 125 481
rect 33 441 125 447
rect 191 481 283 487
rect 191 447 203 481
rect 271 447 283 481
rect 191 441 283 447
rect 349 481 441 487
rect 349 447 361 481
rect 429 447 441 481
rect 349 441 441 447
rect 507 481 599 487
rect 507 447 519 481
rect 587 447 599 481
rect 507 441 599 447
rect 665 481 757 487
rect 665 447 677 481
rect 745 447 757 481
rect 665 441 757 447
rect 823 481 915 487
rect 823 447 835 481
rect 903 447 915 481
rect 823 441 915 447
rect 981 481 1073 487
rect 981 447 993 481
rect 1061 447 1073 481
rect 981 441 1073 447
rect 1139 481 1231 487
rect 1139 447 1151 481
rect 1219 447 1231 481
rect 1139 441 1231 447
rect 1297 481 1389 487
rect 1297 447 1309 481
rect 1377 447 1389 481
rect 1297 441 1389 447
rect 1455 481 1547 487
rect 1455 447 1467 481
rect 1535 447 1547 481
rect 1455 441 1547 447
rect 1613 481 1705 487
rect 1613 447 1625 481
rect 1693 447 1705 481
rect 1613 441 1705 447
rect 1771 481 1863 487
rect 1771 447 1783 481
rect 1851 447 1863 481
rect 1771 441 1863 447
rect 1929 481 2021 487
rect 1929 447 1941 481
rect 2009 447 2021 481
rect 1929 441 2021 447
rect 2087 481 2179 487
rect 2087 447 2099 481
rect 2167 447 2179 481
rect 2087 441 2179 447
rect 2245 481 2337 487
rect 2245 447 2257 481
rect 2325 447 2337 481
rect 2245 441 2337 447
rect 2403 481 2495 487
rect 2403 447 2415 481
rect 2483 447 2495 481
rect 2403 441 2495 447
rect 2561 481 2653 487
rect 2561 447 2573 481
rect 2641 447 2653 481
rect 2561 441 2653 447
rect 2719 481 2811 487
rect 2719 447 2731 481
rect 2799 447 2811 481
rect 2719 441 2811 447
rect 2877 481 2969 487
rect 2877 447 2889 481
rect 2957 447 2969 481
rect 2877 441 2969 447
rect 3035 481 3127 487
rect 3035 447 3047 481
rect 3115 447 3127 481
rect 3035 441 3127 447
rect 3193 481 3285 487
rect 3193 447 3205 481
rect 3273 447 3285 481
rect 3193 441 3285 447
rect 3351 481 3443 487
rect 3351 447 3363 481
rect 3431 447 3443 481
rect 3351 441 3443 447
rect 3509 481 3601 487
rect 3509 447 3521 481
rect 3589 447 3601 481
rect 3509 441 3601 447
rect 3667 481 3759 487
rect 3667 447 3679 481
rect 3747 447 3759 481
rect 3667 441 3759 447
rect 3825 481 3917 487
rect 3825 447 3837 481
rect 3905 447 3917 481
rect 3825 441 3917 447
rect 3983 481 4075 487
rect 3983 447 3995 481
rect 4063 447 4075 481
rect 3983 441 4075 447
rect 4141 481 4233 487
rect 4141 447 4153 481
rect 4221 447 4233 481
rect 4141 441 4233 447
rect 4299 481 4391 487
rect 4299 447 4311 481
rect 4379 447 4391 481
rect 4299 441 4391 447
rect 4457 481 4549 487
rect 4457 447 4469 481
rect 4537 447 4549 481
rect 4457 441 4549 447
rect 4615 481 4707 487
rect 4615 447 4627 481
rect 4695 447 4707 481
rect 4615 441 4707 447
rect 4773 481 4865 487
rect 4773 447 4785 481
rect 4853 447 4865 481
rect 4773 441 4865 447
rect 4931 481 5023 487
rect 4931 447 4943 481
rect 5011 447 5023 481
rect 4931 441 5023 447
rect 5089 481 5181 487
rect 5089 447 5101 481
rect 5169 447 5181 481
rect 5089 441 5181 447
rect 5247 481 5339 487
rect 5247 447 5259 481
rect 5327 447 5339 481
rect 5247 441 5339 447
rect 5405 481 5497 487
rect 5405 447 5417 481
rect 5485 447 5497 481
rect 5405 441 5497 447
rect 5563 481 5655 487
rect 5563 447 5575 481
rect 5643 447 5655 481
rect 5563 441 5655 447
rect 5721 481 5813 487
rect 5721 447 5733 481
rect 5801 447 5813 481
rect 5721 441 5813 447
rect 5879 481 5971 487
rect 5879 447 5891 481
rect 5959 447 5971 481
rect 5879 441 5971 447
rect 6037 481 6129 487
rect 6037 447 6049 481
rect 6117 447 6129 481
rect 6037 441 6129 447
rect 6195 481 6287 487
rect 6195 447 6207 481
rect 6275 447 6287 481
rect 6195 441 6287 447
rect -6343 388 -6297 400
rect -6343 -388 -6337 388
rect -6303 -388 -6297 388
rect -6343 -400 -6297 -388
rect -6185 388 -6139 400
rect -6185 -388 -6179 388
rect -6145 -388 -6139 388
rect -6185 -400 -6139 -388
rect -6027 388 -5981 400
rect -6027 -388 -6021 388
rect -5987 -388 -5981 388
rect -6027 -400 -5981 -388
rect -5869 388 -5823 400
rect -5869 -388 -5863 388
rect -5829 -388 -5823 388
rect -5869 -400 -5823 -388
rect -5711 388 -5665 400
rect -5711 -388 -5705 388
rect -5671 -388 -5665 388
rect -5711 -400 -5665 -388
rect -5553 388 -5507 400
rect -5553 -388 -5547 388
rect -5513 -388 -5507 388
rect -5553 -400 -5507 -388
rect -5395 388 -5349 400
rect -5395 -388 -5389 388
rect -5355 -388 -5349 388
rect -5395 -400 -5349 -388
rect -5237 388 -5191 400
rect -5237 -388 -5231 388
rect -5197 -388 -5191 388
rect -5237 -400 -5191 -388
rect -5079 388 -5033 400
rect -5079 -388 -5073 388
rect -5039 -388 -5033 388
rect -5079 -400 -5033 -388
rect -4921 388 -4875 400
rect -4921 -388 -4915 388
rect -4881 -388 -4875 388
rect -4921 -400 -4875 -388
rect -4763 388 -4717 400
rect -4763 -388 -4757 388
rect -4723 -388 -4717 388
rect -4763 -400 -4717 -388
rect -4605 388 -4559 400
rect -4605 -388 -4599 388
rect -4565 -388 -4559 388
rect -4605 -400 -4559 -388
rect -4447 388 -4401 400
rect -4447 -388 -4441 388
rect -4407 -388 -4401 388
rect -4447 -400 -4401 -388
rect -4289 388 -4243 400
rect -4289 -388 -4283 388
rect -4249 -388 -4243 388
rect -4289 -400 -4243 -388
rect -4131 388 -4085 400
rect -4131 -388 -4125 388
rect -4091 -388 -4085 388
rect -4131 -400 -4085 -388
rect -3973 388 -3927 400
rect -3973 -388 -3967 388
rect -3933 -388 -3927 388
rect -3973 -400 -3927 -388
rect -3815 388 -3769 400
rect -3815 -388 -3809 388
rect -3775 -388 -3769 388
rect -3815 -400 -3769 -388
rect -3657 388 -3611 400
rect -3657 -388 -3651 388
rect -3617 -388 -3611 388
rect -3657 -400 -3611 -388
rect -3499 388 -3453 400
rect -3499 -388 -3493 388
rect -3459 -388 -3453 388
rect -3499 -400 -3453 -388
rect -3341 388 -3295 400
rect -3341 -388 -3335 388
rect -3301 -388 -3295 388
rect -3341 -400 -3295 -388
rect -3183 388 -3137 400
rect -3183 -388 -3177 388
rect -3143 -388 -3137 388
rect -3183 -400 -3137 -388
rect -3025 388 -2979 400
rect -3025 -388 -3019 388
rect -2985 -388 -2979 388
rect -3025 -400 -2979 -388
rect -2867 388 -2821 400
rect -2867 -388 -2861 388
rect -2827 -388 -2821 388
rect -2867 -400 -2821 -388
rect -2709 388 -2663 400
rect -2709 -388 -2703 388
rect -2669 -388 -2663 388
rect -2709 -400 -2663 -388
rect -2551 388 -2505 400
rect -2551 -388 -2545 388
rect -2511 -388 -2505 388
rect -2551 -400 -2505 -388
rect -2393 388 -2347 400
rect -2393 -388 -2387 388
rect -2353 -388 -2347 388
rect -2393 -400 -2347 -388
rect -2235 388 -2189 400
rect -2235 -388 -2229 388
rect -2195 -388 -2189 388
rect -2235 -400 -2189 -388
rect -2077 388 -2031 400
rect -2077 -388 -2071 388
rect -2037 -388 -2031 388
rect -2077 -400 -2031 -388
rect -1919 388 -1873 400
rect -1919 -388 -1913 388
rect -1879 -388 -1873 388
rect -1919 -400 -1873 -388
rect -1761 388 -1715 400
rect -1761 -388 -1755 388
rect -1721 -388 -1715 388
rect -1761 -400 -1715 -388
rect -1603 388 -1557 400
rect -1603 -388 -1597 388
rect -1563 -388 -1557 388
rect -1603 -400 -1557 -388
rect -1445 388 -1399 400
rect -1445 -388 -1439 388
rect -1405 -388 -1399 388
rect -1445 -400 -1399 -388
rect -1287 388 -1241 400
rect -1287 -388 -1281 388
rect -1247 -388 -1241 388
rect -1287 -400 -1241 -388
rect -1129 388 -1083 400
rect -1129 -388 -1123 388
rect -1089 -388 -1083 388
rect -1129 -400 -1083 -388
rect -971 388 -925 400
rect -971 -388 -965 388
rect -931 -388 -925 388
rect -971 -400 -925 -388
rect -813 388 -767 400
rect -813 -388 -807 388
rect -773 -388 -767 388
rect -813 -400 -767 -388
rect -655 388 -609 400
rect -655 -388 -649 388
rect -615 -388 -609 388
rect -655 -400 -609 -388
rect -497 388 -451 400
rect -497 -388 -491 388
rect -457 -388 -451 388
rect -497 -400 -451 -388
rect -339 388 -293 400
rect -339 -388 -333 388
rect -299 -388 -293 388
rect -339 -400 -293 -388
rect -181 388 -135 400
rect -181 -388 -175 388
rect -141 -388 -135 388
rect -181 -400 -135 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 135 388 181 400
rect 135 -388 141 388
rect 175 -388 181 388
rect 135 -400 181 -388
rect 293 388 339 400
rect 293 -388 299 388
rect 333 -388 339 388
rect 293 -400 339 -388
rect 451 388 497 400
rect 451 -388 457 388
rect 491 -388 497 388
rect 451 -400 497 -388
rect 609 388 655 400
rect 609 -388 615 388
rect 649 -388 655 388
rect 609 -400 655 -388
rect 767 388 813 400
rect 767 -388 773 388
rect 807 -388 813 388
rect 767 -400 813 -388
rect 925 388 971 400
rect 925 -388 931 388
rect 965 -388 971 388
rect 925 -400 971 -388
rect 1083 388 1129 400
rect 1083 -388 1089 388
rect 1123 -388 1129 388
rect 1083 -400 1129 -388
rect 1241 388 1287 400
rect 1241 -388 1247 388
rect 1281 -388 1287 388
rect 1241 -400 1287 -388
rect 1399 388 1445 400
rect 1399 -388 1405 388
rect 1439 -388 1445 388
rect 1399 -400 1445 -388
rect 1557 388 1603 400
rect 1557 -388 1563 388
rect 1597 -388 1603 388
rect 1557 -400 1603 -388
rect 1715 388 1761 400
rect 1715 -388 1721 388
rect 1755 -388 1761 388
rect 1715 -400 1761 -388
rect 1873 388 1919 400
rect 1873 -388 1879 388
rect 1913 -388 1919 388
rect 1873 -400 1919 -388
rect 2031 388 2077 400
rect 2031 -388 2037 388
rect 2071 -388 2077 388
rect 2031 -400 2077 -388
rect 2189 388 2235 400
rect 2189 -388 2195 388
rect 2229 -388 2235 388
rect 2189 -400 2235 -388
rect 2347 388 2393 400
rect 2347 -388 2353 388
rect 2387 -388 2393 388
rect 2347 -400 2393 -388
rect 2505 388 2551 400
rect 2505 -388 2511 388
rect 2545 -388 2551 388
rect 2505 -400 2551 -388
rect 2663 388 2709 400
rect 2663 -388 2669 388
rect 2703 -388 2709 388
rect 2663 -400 2709 -388
rect 2821 388 2867 400
rect 2821 -388 2827 388
rect 2861 -388 2867 388
rect 2821 -400 2867 -388
rect 2979 388 3025 400
rect 2979 -388 2985 388
rect 3019 -388 3025 388
rect 2979 -400 3025 -388
rect 3137 388 3183 400
rect 3137 -388 3143 388
rect 3177 -388 3183 388
rect 3137 -400 3183 -388
rect 3295 388 3341 400
rect 3295 -388 3301 388
rect 3335 -388 3341 388
rect 3295 -400 3341 -388
rect 3453 388 3499 400
rect 3453 -388 3459 388
rect 3493 -388 3499 388
rect 3453 -400 3499 -388
rect 3611 388 3657 400
rect 3611 -388 3617 388
rect 3651 -388 3657 388
rect 3611 -400 3657 -388
rect 3769 388 3815 400
rect 3769 -388 3775 388
rect 3809 -388 3815 388
rect 3769 -400 3815 -388
rect 3927 388 3973 400
rect 3927 -388 3933 388
rect 3967 -388 3973 388
rect 3927 -400 3973 -388
rect 4085 388 4131 400
rect 4085 -388 4091 388
rect 4125 -388 4131 388
rect 4085 -400 4131 -388
rect 4243 388 4289 400
rect 4243 -388 4249 388
rect 4283 -388 4289 388
rect 4243 -400 4289 -388
rect 4401 388 4447 400
rect 4401 -388 4407 388
rect 4441 -388 4447 388
rect 4401 -400 4447 -388
rect 4559 388 4605 400
rect 4559 -388 4565 388
rect 4599 -388 4605 388
rect 4559 -400 4605 -388
rect 4717 388 4763 400
rect 4717 -388 4723 388
rect 4757 -388 4763 388
rect 4717 -400 4763 -388
rect 4875 388 4921 400
rect 4875 -388 4881 388
rect 4915 -388 4921 388
rect 4875 -400 4921 -388
rect 5033 388 5079 400
rect 5033 -388 5039 388
rect 5073 -388 5079 388
rect 5033 -400 5079 -388
rect 5191 388 5237 400
rect 5191 -388 5197 388
rect 5231 -388 5237 388
rect 5191 -400 5237 -388
rect 5349 388 5395 400
rect 5349 -388 5355 388
rect 5389 -388 5395 388
rect 5349 -400 5395 -388
rect 5507 388 5553 400
rect 5507 -388 5513 388
rect 5547 -388 5553 388
rect 5507 -400 5553 -388
rect 5665 388 5711 400
rect 5665 -388 5671 388
rect 5705 -388 5711 388
rect 5665 -400 5711 -388
rect 5823 388 5869 400
rect 5823 -388 5829 388
rect 5863 -388 5869 388
rect 5823 -400 5869 -388
rect 5981 388 6027 400
rect 5981 -388 5987 388
rect 6021 -388 6027 388
rect 5981 -400 6027 -388
rect 6139 388 6185 400
rect 6139 -388 6145 388
rect 6179 -388 6185 388
rect 6139 -400 6185 -388
rect 6297 388 6343 400
rect 6297 -388 6303 388
rect 6337 -388 6343 388
rect 6297 -400 6343 -388
rect -6287 -447 -6195 -441
rect -6287 -481 -6275 -447
rect -6207 -481 -6195 -447
rect -6287 -487 -6195 -481
rect -6129 -447 -6037 -441
rect -6129 -481 -6117 -447
rect -6049 -481 -6037 -447
rect -6129 -487 -6037 -481
rect -5971 -447 -5879 -441
rect -5971 -481 -5959 -447
rect -5891 -481 -5879 -447
rect -5971 -487 -5879 -481
rect -5813 -447 -5721 -441
rect -5813 -481 -5801 -447
rect -5733 -481 -5721 -447
rect -5813 -487 -5721 -481
rect -5655 -447 -5563 -441
rect -5655 -481 -5643 -447
rect -5575 -481 -5563 -447
rect -5655 -487 -5563 -481
rect -5497 -447 -5405 -441
rect -5497 -481 -5485 -447
rect -5417 -481 -5405 -447
rect -5497 -487 -5405 -481
rect -5339 -447 -5247 -441
rect -5339 -481 -5327 -447
rect -5259 -481 -5247 -447
rect -5339 -487 -5247 -481
rect -5181 -447 -5089 -441
rect -5181 -481 -5169 -447
rect -5101 -481 -5089 -447
rect -5181 -487 -5089 -481
rect -5023 -447 -4931 -441
rect -5023 -481 -5011 -447
rect -4943 -481 -4931 -447
rect -5023 -487 -4931 -481
rect -4865 -447 -4773 -441
rect -4865 -481 -4853 -447
rect -4785 -481 -4773 -447
rect -4865 -487 -4773 -481
rect -4707 -447 -4615 -441
rect -4707 -481 -4695 -447
rect -4627 -481 -4615 -447
rect -4707 -487 -4615 -481
rect -4549 -447 -4457 -441
rect -4549 -481 -4537 -447
rect -4469 -481 -4457 -447
rect -4549 -487 -4457 -481
rect -4391 -447 -4299 -441
rect -4391 -481 -4379 -447
rect -4311 -481 -4299 -447
rect -4391 -487 -4299 -481
rect -4233 -447 -4141 -441
rect -4233 -481 -4221 -447
rect -4153 -481 -4141 -447
rect -4233 -487 -4141 -481
rect -4075 -447 -3983 -441
rect -4075 -481 -4063 -447
rect -3995 -481 -3983 -447
rect -4075 -487 -3983 -481
rect -3917 -447 -3825 -441
rect -3917 -481 -3905 -447
rect -3837 -481 -3825 -447
rect -3917 -487 -3825 -481
rect -3759 -447 -3667 -441
rect -3759 -481 -3747 -447
rect -3679 -481 -3667 -447
rect -3759 -487 -3667 -481
rect -3601 -447 -3509 -441
rect -3601 -481 -3589 -447
rect -3521 -481 -3509 -447
rect -3601 -487 -3509 -481
rect -3443 -447 -3351 -441
rect -3443 -481 -3431 -447
rect -3363 -481 -3351 -447
rect -3443 -487 -3351 -481
rect -3285 -447 -3193 -441
rect -3285 -481 -3273 -447
rect -3205 -481 -3193 -447
rect -3285 -487 -3193 -481
rect -3127 -447 -3035 -441
rect -3127 -481 -3115 -447
rect -3047 -481 -3035 -447
rect -3127 -487 -3035 -481
rect -2969 -447 -2877 -441
rect -2969 -481 -2957 -447
rect -2889 -481 -2877 -447
rect -2969 -487 -2877 -481
rect -2811 -447 -2719 -441
rect -2811 -481 -2799 -447
rect -2731 -481 -2719 -447
rect -2811 -487 -2719 -481
rect -2653 -447 -2561 -441
rect -2653 -481 -2641 -447
rect -2573 -481 -2561 -447
rect -2653 -487 -2561 -481
rect -2495 -447 -2403 -441
rect -2495 -481 -2483 -447
rect -2415 -481 -2403 -447
rect -2495 -487 -2403 -481
rect -2337 -447 -2245 -441
rect -2337 -481 -2325 -447
rect -2257 -481 -2245 -447
rect -2337 -487 -2245 -481
rect -2179 -447 -2087 -441
rect -2179 -481 -2167 -447
rect -2099 -481 -2087 -447
rect -2179 -487 -2087 -481
rect -2021 -447 -1929 -441
rect -2021 -481 -2009 -447
rect -1941 -481 -1929 -447
rect -2021 -487 -1929 -481
rect -1863 -447 -1771 -441
rect -1863 -481 -1851 -447
rect -1783 -481 -1771 -447
rect -1863 -487 -1771 -481
rect -1705 -447 -1613 -441
rect -1705 -481 -1693 -447
rect -1625 -481 -1613 -447
rect -1705 -487 -1613 -481
rect -1547 -447 -1455 -441
rect -1547 -481 -1535 -447
rect -1467 -481 -1455 -447
rect -1547 -487 -1455 -481
rect -1389 -447 -1297 -441
rect -1389 -481 -1377 -447
rect -1309 -481 -1297 -447
rect -1389 -487 -1297 -481
rect -1231 -447 -1139 -441
rect -1231 -481 -1219 -447
rect -1151 -481 -1139 -447
rect -1231 -487 -1139 -481
rect -1073 -447 -981 -441
rect -1073 -481 -1061 -447
rect -993 -481 -981 -447
rect -1073 -487 -981 -481
rect -915 -447 -823 -441
rect -915 -481 -903 -447
rect -835 -481 -823 -447
rect -915 -487 -823 -481
rect -757 -447 -665 -441
rect -757 -481 -745 -447
rect -677 -481 -665 -447
rect -757 -487 -665 -481
rect -599 -447 -507 -441
rect -599 -481 -587 -447
rect -519 -481 -507 -447
rect -599 -487 -507 -481
rect -441 -447 -349 -441
rect -441 -481 -429 -447
rect -361 -481 -349 -447
rect -441 -487 -349 -481
rect -283 -447 -191 -441
rect -283 -481 -271 -447
rect -203 -481 -191 -447
rect -283 -487 -191 -481
rect -125 -447 -33 -441
rect -125 -481 -113 -447
rect -45 -481 -33 -447
rect -125 -487 -33 -481
rect 33 -447 125 -441
rect 33 -481 45 -447
rect 113 -481 125 -447
rect 33 -487 125 -481
rect 191 -447 283 -441
rect 191 -481 203 -447
rect 271 -481 283 -447
rect 191 -487 283 -481
rect 349 -447 441 -441
rect 349 -481 361 -447
rect 429 -481 441 -447
rect 349 -487 441 -481
rect 507 -447 599 -441
rect 507 -481 519 -447
rect 587 -481 599 -447
rect 507 -487 599 -481
rect 665 -447 757 -441
rect 665 -481 677 -447
rect 745 -481 757 -447
rect 665 -487 757 -481
rect 823 -447 915 -441
rect 823 -481 835 -447
rect 903 -481 915 -447
rect 823 -487 915 -481
rect 981 -447 1073 -441
rect 981 -481 993 -447
rect 1061 -481 1073 -447
rect 981 -487 1073 -481
rect 1139 -447 1231 -441
rect 1139 -481 1151 -447
rect 1219 -481 1231 -447
rect 1139 -487 1231 -481
rect 1297 -447 1389 -441
rect 1297 -481 1309 -447
rect 1377 -481 1389 -447
rect 1297 -487 1389 -481
rect 1455 -447 1547 -441
rect 1455 -481 1467 -447
rect 1535 -481 1547 -447
rect 1455 -487 1547 -481
rect 1613 -447 1705 -441
rect 1613 -481 1625 -447
rect 1693 -481 1705 -447
rect 1613 -487 1705 -481
rect 1771 -447 1863 -441
rect 1771 -481 1783 -447
rect 1851 -481 1863 -447
rect 1771 -487 1863 -481
rect 1929 -447 2021 -441
rect 1929 -481 1941 -447
rect 2009 -481 2021 -447
rect 1929 -487 2021 -481
rect 2087 -447 2179 -441
rect 2087 -481 2099 -447
rect 2167 -481 2179 -447
rect 2087 -487 2179 -481
rect 2245 -447 2337 -441
rect 2245 -481 2257 -447
rect 2325 -481 2337 -447
rect 2245 -487 2337 -481
rect 2403 -447 2495 -441
rect 2403 -481 2415 -447
rect 2483 -481 2495 -447
rect 2403 -487 2495 -481
rect 2561 -447 2653 -441
rect 2561 -481 2573 -447
rect 2641 -481 2653 -447
rect 2561 -487 2653 -481
rect 2719 -447 2811 -441
rect 2719 -481 2731 -447
rect 2799 -481 2811 -447
rect 2719 -487 2811 -481
rect 2877 -447 2969 -441
rect 2877 -481 2889 -447
rect 2957 -481 2969 -447
rect 2877 -487 2969 -481
rect 3035 -447 3127 -441
rect 3035 -481 3047 -447
rect 3115 -481 3127 -447
rect 3035 -487 3127 -481
rect 3193 -447 3285 -441
rect 3193 -481 3205 -447
rect 3273 -481 3285 -447
rect 3193 -487 3285 -481
rect 3351 -447 3443 -441
rect 3351 -481 3363 -447
rect 3431 -481 3443 -447
rect 3351 -487 3443 -481
rect 3509 -447 3601 -441
rect 3509 -481 3521 -447
rect 3589 -481 3601 -447
rect 3509 -487 3601 -481
rect 3667 -447 3759 -441
rect 3667 -481 3679 -447
rect 3747 -481 3759 -447
rect 3667 -487 3759 -481
rect 3825 -447 3917 -441
rect 3825 -481 3837 -447
rect 3905 -481 3917 -447
rect 3825 -487 3917 -481
rect 3983 -447 4075 -441
rect 3983 -481 3995 -447
rect 4063 -481 4075 -447
rect 3983 -487 4075 -481
rect 4141 -447 4233 -441
rect 4141 -481 4153 -447
rect 4221 -481 4233 -447
rect 4141 -487 4233 -481
rect 4299 -447 4391 -441
rect 4299 -481 4311 -447
rect 4379 -481 4391 -447
rect 4299 -487 4391 -481
rect 4457 -447 4549 -441
rect 4457 -481 4469 -447
rect 4537 -481 4549 -447
rect 4457 -487 4549 -481
rect 4615 -447 4707 -441
rect 4615 -481 4627 -447
rect 4695 -481 4707 -447
rect 4615 -487 4707 -481
rect 4773 -447 4865 -441
rect 4773 -481 4785 -447
rect 4853 -481 4865 -447
rect 4773 -487 4865 -481
rect 4931 -447 5023 -441
rect 4931 -481 4943 -447
rect 5011 -481 5023 -447
rect 4931 -487 5023 -481
rect 5089 -447 5181 -441
rect 5089 -481 5101 -447
rect 5169 -481 5181 -447
rect 5089 -487 5181 -481
rect 5247 -447 5339 -441
rect 5247 -481 5259 -447
rect 5327 -481 5339 -447
rect 5247 -487 5339 -481
rect 5405 -447 5497 -441
rect 5405 -481 5417 -447
rect 5485 -481 5497 -447
rect 5405 -487 5497 -481
rect 5563 -447 5655 -441
rect 5563 -481 5575 -447
rect 5643 -481 5655 -447
rect 5563 -487 5655 -481
rect 5721 -447 5813 -441
rect 5721 -481 5733 -447
rect 5801 -481 5813 -447
rect 5721 -487 5813 -481
rect 5879 -447 5971 -441
rect 5879 -481 5891 -447
rect 5959 -481 5971 -447
rect 5879 -487 5971 -481
rect 6037 -447 6129 -441
rect 6037 -481 6049 -447
rect 6117 -481 6129 -447
rect 6037 -487 6129 -481
rect 6195 -447 6287 -441
rect 6195 -481 6207 -447
rect 6275 -481 6287 -447
rect 6195 -487 6287 -481
<< properties >>
string FIXED_BBOX -6454 -602 6454 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.50 m 1 nf 80 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
