magic
tech sky130A
timestamp 1666553597
<< metal4 >>
rect -10078 1679 -6825 3125
rect -6785 1679 -3532 3125
rect -3492 1679 -221 3125
rect -181 1679 3090 3125
rect 3130 1679 6384 3125
rect 6424 1679 9778 3125
rect -10078 1490 9778 1679
rect -10078 25 -6825 1490
rect -6785 25 -3532 1490
rect -3492 25 -221 1490
rect -181 25 3090 1490
rect 3130 25 6384 1490
rect 6424 25 9778 1490
rect -8608 -25 -8447 25
rect -5316 -25 -5155 25
rect -2023 -25 -1862 25
rect 1288 -25 1449 25
rect 4600 -25 4761 25
rect 7897 -25 8058 25
rect -10078 -1516 -6825 -25
rect -6785 -1516 -3532 -25
rect -3492 -1516 -221 -25
rect -181 -1516 3090 -25
rect 3130 -1516 6384 -25
rect 6424 -1516 9778 -25
rect -10078 -1705 9778 -1516
rect -10078 -3125 -6825 -1705
rect -6785 -3125 -3532 -1705
rect -3492 -3125 -221 -1705
rect -181 -3125 3090 -1705
rect 3130 -3125 6384 -1705
rect 6424 -3125 9778 -1705
<< mimcap2 >>
rect -10028 3055 -7028 3075
rect -10028 95 -10008 3055
rect -7048 95 -7028 3055
rect -10028 75 -7028 95
rect -6735 3055 -3735 3075
rect -6735 95 -6715 3055
rect -3755 95 -3735 3055
rect -6735 75 -3735 95
rect -3442 3055 -442 3075
rect -3442 95 -3422 3055
rect -462 95 -442 3055
rect -3442 75 -442 95
rect -131 3055 2869 3075
rect -131 95 -111 3055
rect 2849 95 2869 3055
rect -131 75 2869 95
rect 3180 3055 6180 3075
rect 3180 95 3200 3055
rect 6160 95 6180 3055
rect 3180 75 6180 95
rect 6474 3055 9477 3075
rect 6474 95 6494 3055
rect 9457 95 9477 3055
rect 6474 75 9477 95
rect -10028 -95 -7028 -75
rect -10028 -3055 -10008 -95
rect -7048 -3055 -7028 -95
rect -10028 -3075 -7028 -3055
rect -6735 -95 -3735 -75
rect -6735 -3055 -6715 -95
rect -3755 -3055 -3735 -95
rect -6735 -3075 -3735 -3055
rect -3442 -95 -442 -75
rect -3442 -3055 -3422 -95
rect -462 -3055 -442 -95
rect -3442 -3075 -442 -3055
rect -131 -95 2869 -75
rect -131 -3055 -111 -95
rect 2849 -3055 2869 -95
rect -131 -3075 2869 -3055
rect 3180 -95 6180 -75
rect 3180 -3055 3200 -95
rect 6160 -3055 6180 -95
rect 3180 -3075 6180 -3055
rect 6474 -95 9477 -75
rect 6474 -3055 6494 -95
rect 9457 -3055 9477 -95
rect 6474 -3075 9477 -3055
<< mimcap2contact >>
rect -10008 95 -7048 3055
rect -6715 95 -3755 3055
rect -3422 95 -462 3055
rect -111 95 2849 3055
rect 3200 95 6160 3055
rect 6494 95 9457 3055
rect -10008 -3055 -7048 -95
rect -6715 -3055 -3755 -95
rect -3422 -3055 -462 -95
rect -111 -3055 2849 -95
rect 3200 -3055 6160 -95
rect 6494 -3055 9457 -95
<< metal5 >>
rect -8608 3067 -8448 3150
rect -7048 3067 -6888 3150
rect -5315 3067 -5155 3150
rect -3755 3067 -3595 3150
rect -2022 3067 -1862 3150
rect -462 3067 -302 3150
rect 1289 3067 1449 3150
rect 2849 3067 3009 3150
rect 4600 3067 4760 3150
rect 6160 3067 6320 3150
rect 7897 3067 8057 3150
rect 9457 3067 9617 3150
rect -10020 3055 -6888 3067
rect -10020 95 -10008 3055
rect -7048 1679 -6888 3055
rect -6727 3055 -3595 3067
rect -6727 1679 -6715 3055
rect -7048 1490 -6715 1679
rect -7048 95 -6888 1490
rect -10020 83 -6888 95
rect -6727 95 -6715 1490
rect -3755 1679 -3595 3055
rect -3434 3055 -302 3067
rect -3434 1679 -3422 3055
rect -3755 1490 -3422 1679
rect -3755 95 -3595 1490
rect -6727 83 -3595 95
rect -3434 95 -3422 1490
rect -462 1679 -302 3055
rect -123 3055 3009 3067
rect -123 1679 -111 3055
rect -462 1490 -111 1679
rect -462 95 -302 1490
rect -3434 83 -302 95
rect -123 95 -111 1490
rect 2849 1679 3009 3055
rect 3188 3055 6320 3067
rect 3188 1679 3200 3055
rect 2849 1490 3200 1679
rect 2849 95 3009 1490
rect -123 83 3009 95
rect 3188 95 3200 1490
rect 6160 1679 6320 3055
rect 6482 3055 9617 3067
rect 6482 1679 6494 3055
rect 6160 1490 6494 1679
rect 6160 95 6320 1490
rect 3188 83 6320 95
rect 6482 95 6494 1490
rect 9457 95 9617 3055
rect 6482 83 9617 95
rect -8608 -83 -8448 83
rect -7048 -83 -6888 83
rect -5315 -83 -5155 83
rect -3755 -83 -3595 83
rect -2022 -83 -1862 83
rect -462 -83 -302 83
rect 1289 -83 1449 83
rect 2849 -83 3009 83
rect 4600 -83 4760 83
rect 6160 -83 6320 83
rect 7897 -83 8057 83
rect 9457 -83 9617 83
rect -10020 -95 -6888 -83
rect -10020 -3055 -10008 -95
rect -7048 -1516 -6888 -95
rect -6727 -95 -3595 -83
rect -6727 -1516 -6715 -95
rect -7048 -1705 -6715 -1516
rect -7048 -3055 -6888 -1705
rect -10020 -3067 -6888 -3055
rect -6727 -3055 -6715 -1705
rect -3755 -1516 -3595 -95
rect -3434 -95 -302 -83
rect -3434 -1516 -3422 -95
rect -3755 -1705 -3422 -1516
rect -3755 -3055 -3595 -1705
rect -6727 -3067 -3595 -3055
rect -3434 -3055 -3422 -1705
rect -462 -1516 -302 -95
rect -123 -95 3009 -83
rect -123 -1516 -111 -95
rect -462 -1705 -111 -1516
rect -462 -3055 -302 -1705
rect -3434 -3067 -302 -3055
rect -123 -3055 -111 -1705
rect 2849 -1516 3009 -95
rect 3188 -95 6320 -83
rect 3188 -1516 3200 -95
rect 2849 -1705 3200 -1516
rect 2849 -3055 3009 -1705
rect -123 -3067 3009 -3055
rect 3188 -3055 3200 -1705
rect 6160 -1516 6320 -95
rect 6482 -95 9617 -83
rect 6482 -1516 6494 -95
rect 6160 -1705 6494 -1516
rect 6160 -3055 6320 -1705
rect 3188 -3067 6320 -3055
rect 6482 -3055 6494 -1705
rect 9457 -3055 9617 -95
rect 6482 -3067 9617 -3055
rect -8608 -3150 -8448 -3067
rect -7048 -3150 -6888 -3067
rect -5315 -3150 -5155 -3067
rect -3755 -3150 -3595 -3067
rect -2022 -3150 -1862 -3067
rect -462 -3150 -302 -3067
rect 1289 -3150 1449 -3067
rect 2849 -3150 3009 -3067
rect 4600 -3150 4760 -3067
rect 6160 -3150 6320 -3067
rect 7897 -3150 8057 -3067
rect 9457 -3150 9617 -3067
<< properties >>
string FIXED_BBOX 6727 25 9827 3125
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 6 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
