magic
tech sky130A
magscale 1 2
timestamp 1666207736
<< error_p >>
rect -2895 2865 -2835 8395
rect -2815 2865 -2755 8395
rect 2754 2865 2814 8395
rect 2834 2865 2894 8395
rect -2895 -2765 -2835 2765
rect -2815 -2765 -2755 2765
rect 2754 -2765 2814 2765
rect 2834 -2765 2894 2765
rect -2895 -8395 -2835 -2865
rect -2815 -8395 -2755 -2865
rect 2754 -8395 2814 -2865
rect 2834 -8395 2894 -2865
<< metal3 >>
rect -8464 8367 -2835 8395
rect -8464 2893 -2919 8367
rect -2855 2893 -2835 8367
rect -8464 2865 -2835 2893
rect -2815 8367 2814 8395
rect -2815 2893 2730 8367
rect 2794 2893 2814 8367
rect -2815 2865 2814 2893
rect 2834 8367 8463 8395
rect 2834 2893 8379 8367
rect 8443 2893 8463 8367
rect 2834 2865 8463 2893
rect -8464 2737 -2835 2765
rect -8464 -2737 -2919 2737
rect -2855 -2737 -2835 2737
rect -8464 -2765 -2835 -2737
rect -2815 2737 2814 2765
rect -2815 -2737 2730 2737
rect 2794 -2737 2814 2737
rect -2815 -2765 2814 -2737
rect 2834 2737 8463 2765
rect 2834 -2737 8379 2737
rect 8443 -2737 8463 2737
rect 2834 -2765 8463 -2737
rect -8464 -2893 -2835 -2865
rect -8464 -8367 -2919 -2893
rect -2855 -8367 -2835 -2893
rect -8464 -8395 -2835 -8367
rect -2815 -2893 2814 -2865
rect -2815 -8367 2730 -2893
rect 2794 -8367 2814 -2893
rect -2815 -8395 2814 -8367
rect 2834 -2893 8463 -2865
rect 2834 -8367 8379 -2893
rect 8443 -8367 8463 -2893
rect 2834 -8395 8463 -8367
<< via3 >>
rect -2919 2893 -2855 8367
rect 2730 2893 2794 8367
rect 8379 2893 8443 8367
rect -2919 -2737 -2855 2737
rect 2730 -2737 2794 2737
rect 8379 -2737 8443 2737
rect -2919 -8367 -2855 -2893
rect 2730 -8367 2794 -2893
rect 8379 -8367 8443 -2893
<< mimcap >>
rect -8364 8255 -3034 8295
rect -8364 3005 -8324 8255
rect -3074 3005 -3034 8255
rect -8364 2965 -3034 3005
rect -2715 8255 2615 8295
rect -2715 3005 -2675 8255
rect 2575 3005 2615 8255
rect -2715 2965 2615 3005
rect 2934 8255 8264 8295
rect 2934 3005 2974 8255
rect 8224 3005 8264 8255
rect 2934 2965 8264 3005
rect -8364 2625 -3034 2665
rect -8364 -2625 -8324 2625
rect -3074 -2625 -3034 2625
rect -8364 -2665 -3034 -2625
rect -2715 2625 2615 2665
rect -2715 -2625 -2675 2625
rect 2575 -2625 2615 2625
rect -2715 -2665 2615 -2625
rect 2934 2625 8264 2665
rect 2934 -2625 2974 2625
rect 8224 -2625 8264 2625
rect 2934 -2665 8264 -2625
rect -8364 -3005 -3034 -2965
rect -8364 -8255 -8324 -3005
rect -3074 -8255 -3034 -3005
rect -8364 -8295 -3034 -8255
rect -2715 -3005 2615 -2965
rect -2715 -8255 -2675 -3005
rect 2575 -8255 2615 -3005
rect -2715 -8295 2615 -8255
rect 2934 -3005 8264 -2965
rect 2934 -8255 2974 -3005
rect 8224 -8255 8264 -3005
rect 2934 -8295 8264 -8255
<< mimcapcontact >>
rect -8324 3005 -3074 8255
rect -2675 3005 2575 8255
rect 2974 3005 8224 8255
rect -8324 -2625 -3074 2625
rect -2675 -2625 2575 2625
rect 2974 -2625 8224 2625
rect -8324 -8255 -3074 -3005
rect -2675 -8255 2575 -3005
rect 2974 -8255 8224 -3005
<< metal4 >>
rect -5751 8256 -5647 8445
rect -2966 8383 -2862 8445
rect -2966 8367 -2839 8383
rect -8325 8255 -3073 8256
rect -8325 3005 -8324 8255
rect -3074 3005 -3073 8255
rect -8325 3004 -3073 3005
rect -5751 2626 -5647 3004
rect -2966 2893 -2919 8367
rect -2855 2893 -2839 8367
rect -102 8256 2 8445
rect 2683 8383 2787 8445
rect 2683 8367 2810 8383
rect -2676 8255 2576 8256
rect -2676 3005 -2675 8255
rect 2575 3005 2576 8255
rect -2676 3004 2576 3005
rect -2966 2877 -2839 2893
rect -2966 2753 -2862 2877
rect -2966 2737 -2839 2753
rect -8325 2625 -3073 2626
rect -8325 -2625 -8324 2625
rect -3074 -2625 -3073 2625
rect -8325 -2626 -3073 -2625
rect -5751 -3004 -5647 -2626
rect -2966 -2737 -2919 2737
rect -2855 -2737 -2839 2737
rect -102 2626 2 3004
rect 2683 2893 2730 8367
rect 2794 2893 2810 8367
rect 5547 8256 5651 8445
rect 8332 8383 8436 8445
rect 8332 8367 8459 8383
rect 2973 8255 8225 8256
rect 2973 3005 2974 8255
rect 8224 3005 8225 8255
rect 2973 3004 8225 3005
rect 2683 2877 2810 2893
rect 2683 2753 2787 2877
rect 2683 2737 2810 2753
rect -2676 2625 2576 2626
rect -2676 -2625 -2675 2625
rect 2575 -2625 2576 2625
rect -2676 -2626 2576 -2625
rect -2966 -2753 -2839 -2737
rect -2966 -2877 -2862 -2753
rect -2966 -2893 -2839 -2877
rect -8325 -3005 -3073 -3004
rect -8325 -8255 -8324 -3005
rect -3074 -8255 -3073 -3005
rect -8325 -8256 -3073 -8255
rect -5751 -8445 -5647 -8256
rect -2966 -8367 -2919 -2893
rect -2855 -8367 -2839 -2893
rect -102 -3004 2 -2626
rect 2683 -2737 2730 2737
rect 2794 -2737 2810 2737
rect 5547 2626 5651 3004
rect 8332 2893 8379 8367
rect 8443 2893 8459 8367
rect 8332 2877 8459 2893
rect 8332 2753 8436 2877
rect 8332 2737 8459 2753
rect 2973 2625 8225 2626
rect 2973 -2625 2974 2625
rect 8224 -2625 8225 2625
rect 2973 -2626 8225 -2625
rect 2683 -2753 2810 -2737
rect 2683 -2877 2787 -2753
rect 2683 -2893 2810 -2877
rect -2676 -3005 2576 -3004
rect -2676 -8255 -2675 -3005
rect 2575 -8255 2576 -3005
rect -2676 -8256 2576 -8255
rect -2966 -8383 -2839 -8367
rect -2966 -8445 -2862 -8383
rect -102 -8445 2 -8256
rect 2683 -8367 2730 -2893
rect 2794 -8367 2810 -2893
rect 5547 -3004 5651 -2626
rect 8332 -2737 8379 2737
rect 8443 -2737 8459 2737
rect 8332 -2753 8459 -2737
rect 8332 -2877 8436 -2753
rect 8332 -2893 8459 -2877
rect 2973 -3005 8225 -3004
rect 2973 -8255 2974 -3005
rect 8224 -8255 8225 -3005
rect 2973 -8256 8225 -8255
rect 2683 -8383 2810 -8367
rect 2683 -8445 2787 -8383
rect 5547 -8445 5651 -8256
rect 8332 -8367 8379 -2893
rect 8443 -8367 8459 -2893
rect 8332 -8383 8459 -8367
rect 8332 -8445 8436 -8383
<< properties >>
string FIXED_BBOX 2834 2865 8364 8395
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 26.65 l 26.65 val 1.44k carea 2.00 cperi 0.19 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
