magic
tech sky130A
magscale 1 2
timestamp 1668293870
<< pwell >>
rect -783 -710 783 710
<< nmos >>
rect -587 -500 -337 500
rect -279 -500 -29 500
rect 29 -500 279 500
rect 337 -500 587 500
<< ndiff >>
rect -645 488 -587 500
rect -645 -488 -633 488
rect -599 -488 -587 488
rect -645 -500 -587 -488
rect -337 488 -279 500
rect -337 -488 -325 488
rect -291 -488 -279 488
rect -337 -500 -279 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 279 488 337 500
rect 279 -488 291 488
rect 325 -488 337 488
rect 279 -500 337 -488
rect 587 488 645 500
rect 587 -488 599 488
rect 633 -488 645 488
rect 587 -500 645 -488
<< ndiffc >>
rect -633 -488 -599 488
rect -325 -488 -291 488
rect -17 -488 17 488
rect 291 -488 325 488
rect 599 -488 633 488
<< psubdiff >>
rect -747 640 -651 674
rect 651 640 747 674
rect -747 578 -713 640
rect 713 578 747 640
rect -747 -640 -713 -578
rect 713 -640 747 -578
rect -747 -674 -651 -640
rect 651 -674 747 -640
<< psubdiffcont >>
rect -651 640 651 674
rect -747 -578 -713 578
rect 713 -578 747 578
rect -651 -674 651 -640
<< poly >>
rect -587 572 -337 588
rect -587 538 -571 572
rect -353 538 -337 572
rect -587 500 -337 538
rect -279 572 -29 588
rect -279 538 -263 572
rect -45 538 -29 572
rect -279 500 -29 538
rect 29 572 279 588
rect 29 538 45 572
rect 263 538 279 572
rect 29 500 279 538
rect 337 572 587 588
rect 337 538 353 572
rect 571 538 587 572
rect 337 500 587 538
rect -587 -538 -337 -500
rect -587 -572 -571 -538
rect -353 -572 -337 -538
rect -587 -588 -337 -572
rect -279 -538 -29 -500
rect -279 -572 -263 -538
rect -45 -572 -29 -538
rect -279 -588 -29 -572
rect 29 -538 279 -500
rect 29 -572 45 -538
rect 263 -572 279 -538
rect 29 -588 279 -572
rect 337 -538 587 -500
rect 337 -572 353 -538
rect 571 -572 587 -538
rect 337 -588 587 -572
<< polycont >>
rect -571 538 -353 572
rect -263 538 -45 572
rect 45 538 263 572
rect 353 538 571 572
rect -571 -572 -353 -538
rect -263 -572 -45 -538
rect 45 -572 263 -538
rect 353 -572 571 -538
<< locali >>
rect -747 640 -651 674
rect 651 640 747 674
rect -747 578 -713 640
rect 713 578 747 640
rect -587 538 -571 572
rect -353 538 -337 572
rect -279 538 -263 572
rect -45 538 -29 572
rect 29 538 45 572
rect 263 538 279 572
rect 337 538 353 572
rect 571 538 587 572
rect -633 488 -599 504
rect -633 -504 -599 -488
rect -325 488 -291 504
rect -325 -504 -291 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 291 488 325 504
rect 291 -504 325 -488
rect 599 488 633 504
rect 599 -504 633 -488
rect -587 -572 -571 -538
rect -353 -572 -337 -538
rect -279 -572 -263 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 263 -572 279 -538
rect 337 -572 353 -538
rect 571 -572 587 -538
rect -747 -640 -713 -578
rect 713 -640 747 -578
rect -747 -674 -651 -640
rect 651 -674 747 -640
<< viali >>
rect -571 538 -353 572
rect -263 538 -45 572
rect 45 538 263 572
rect 353 538 571 572
rect -633 -488 -599 488
rect -325 -488 -291 488
rect -17 -488 17 488
rect 291 -488 325 488
rect 599 -488 633 488
rect -571 -572 -353 -538
rect -263 -572 -45 -538
rect 45 -572 263 -538
rect 353 -572 571 -538
<< metal1 >>
rect -583 572 -341 578
rect -583 538 -571 572
rect -353 538 -341 572
rect -583 532 -341 538
rect -275 572 -33 578
rect -275 538 -263 572
rect -45 538 -33 572
rect -275 532 -33 538
rect 33 572 275 578
rect 33 538 45 572
rect 263 538 275 572
rect 33 532 275 538
rect 341 572 583 578
rect 341 538 353 572
rect 571 538 583 572
rect 341 532 583 538
rect -639 488 -593 500
rect -639 -488 -633 488
rect -599 -488 -593 488
rect -639 -500 -593 -488
rect -331 488 -285 500
rect -331 -488 -325 488
rect -291 -488 -285 488
rect -331 -500 -285 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 285 488 331 500
rect 285 -488 291 488
rect 325 -488 331 488
rect 285 -500 331 -488
rect 593 488 639 500
rect 593 -488 599 488
rect 633 -488 639 488
rect 593 -500 639 -488
rect -583 -538 -341 -532
rect -583 -572 -571 -538
rect -353 -572 -341 -538
rect -583 -578 -341 -572
rect -275 -538 -33 -532
rect -275 -572 -263 -538
rect -45 -572 -33 -538
rect -275 -578 -33 -572
rect 33 -538 275 -532
rect 33 -572 45 -538
rect 263 -572 275 -538
rect 33 -578 275 -572
rect 341 -538 583 -532
rect 341 -572 353 -538
rect 571 -572 583 -538
rect 341 -578 583 -572
<< properties >>
string FIXED_BBOX -730 -657 730 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
