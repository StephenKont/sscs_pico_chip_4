magic
tech sky130A
timestamp 1667069478
<< pwell >>
rect -1422 -1129 1422 1129
<< mvnmos >>
rect -1308 -1000 -808 1000
rect -779 -1000 -279 1000
rect -250 -1000 250 1000
rect 279 -1000 779 1000
rect 808 -1000 1308 1000
<< mvndiff >>
rect -1337 994 -1308 1000
rect -1337 -994 -1331 994
rect -1314 -994 -1308 994
rect -1337 -1000 -1308 -994
rect -808 994 -779 1000
rect -808 -994 -802 994
rect -785 -994 -779 994
rect -808 -1000 -779 -994
rect -279 994 -250 1000
rect -279 -994 -273 994
rect -256 -994 -250 994
rect -279 -1000 -250 -994
rect 250 994 279 1000
rect 250 -994 256 994
rect 273 -994 279 994
rect 250 -1000 279 -994
rect 779 994 808 1000
rect 779 -994 785 994
rect 802 -994 808 994
rect 779 -1000 808 -994
rect 1308 994 1337 1000
rect 1308 -994 1314 994
rect 1331 -994 1337 994
rect 1308 -1000 1337 -994
<< mvndiffc >>
rect -1331 -994 -1314 994
rect -802 -994 -785 994
rect -273 -994 -256 994
rect 256 -994 273 994
rect 785 -994 802 994
rect 1314 -994 1331 994
<< mvpsubdiff >>
rect -1404 1105 1404 1111
rect -1404 1088 -1350 1105
rect 1350 1088 1404 1105
rect -1404 1082 1404 1088
rect -1404 1057 -1375 1082
rect -1404 -1057 -1398 1057
rect -1381 -1057 -1375 1057
rect 1375 1057 1404 1082
rect -1404 -1082 -1375 -1057
rect 1375 -1057 1381 1057
rect 1398 -1057 1404 1057
rect 1375 -1082 1404 -1057
rect -1404 -1088 1404 -1082
rect -1404 -1105 -1350 -1088
rect 1350 -1105 1404 -1088
rect -1404 -1111 1404 -1105
<< mvpsubdiffcont >>
rect -1350 1088 1350 1105
rect -1398 -1057 -1381 1057
rect 1381 -1057 1398 1057
rect -1350 -1105 1350 -1088
<< poly >>
rect -1308 1036 -808 1044
rect -1308 1019 -1300 1036
rect -816 1019 -808 1036
rect -1308 1000 -808 1019
rect -779 1036 -279 1044
rect -779 1019 -771 1036
rect -287 1019 -279 1036
rect -779 1000 -279 1019
rect -250 1036 250 1044
rect -250 1019 -242 1036
rect 242 1019 250 1036
rect -250 1000 250 1019
rect 279 1036 779 1044
rect 279 1019 287 1036
rect 771 1019 779 1036
rect 279 1000 779 1019
rect 808 1036 1308 1044
rect 808 1019 816 1036
rect 1300 1019 1308 1036
rect 808 1000 1308 1019
rect -1308 -1019 -808 -1000
rect -1308 -1036 -1300 -1019
rect -816 -1036 -808 -1019
rect -1308 -1044 -808 -1036
rect -779 -1019 -279 -1000
rect -779 -1036 -771 -1019
rect -287 -1036 -279 -1019
rect -779 -1044 -279 -1036
rect -250 -1019 250 -1000
rect -250 -1036 -242 -1019
rect 242 -1036 250 -1019
rect -250 -1044 250 -1036
rect 279 -1019 779 -1000
rect 279 -1036 287 -1019
rect 771 -1036 779 -1019
rect 279 -1044 779 -1036
rect 808 -1019 1308 -1000
rect 808 -1036 816 -1019
rect 1300 -1036 1308 -1019
rect 808 -1044 1308 -1036
<< polycont >>
rect -1300 1019 -816 1036
rect -771 1019 -287 1036
rect -242 1019 242 1036
rect 287 1019 771 1036
rect 816 1019 1300 1036
rect -1300 -1036 -816 -1019
rect -771 -1036 -287 -1019
rect -242 -1036 242 -1019
rect 287 -1036 771 -1019
rect 816 -1036 1300 -1019
<< locali >>
rect -1398 1088 -1350 1105
rect 1350 1088 1398 1105
rect -1398 1057 -1381 1088
rect 1381 1057 1398 1088
rect -1308 1019 -1300 1036
rect -816 1019 -808 1036
rect -779 1019 -771 1036
rect -287 1019 -279 1036
rect -250 1019 -242 1036
rect 242 1019 250 1036
rect 279 1019 287 1036
rect 771 1019 779 1036
rect 808 1019 816 1036
rect 1300 1019 1308 1036
rect -1331 994 -1314 1002
rect -1331 -1002 -1314 -994
rect -802 994 -785 1002
rect -802 -1002 -785 -994
rect -273 994 -256 1002
rect -273 -1002 -256 -994
rect 256 994 273 1002
rect 256 -1002 273 -994
rect 785 994 802 1002
rect 785 -1002 802 -994
rect 1314 994 1331 1002
rect 1314 -1002 1331 -994
rect -1308 -1036 -1300 -1019
rect -816 -1036 -808 -1019
rect -779 -1036 -771 -1019
rect -287 -1036 -279 -1019
rect -250 -1036 -242 -1019
rect 242 -1036 250 -1019
rect 279 -1036 287 -1019
rect 771 -1036 779 -1019
rect 808 -1036 816 -1019
rect 1300 -1036 1308 -1019
rect -1398 -1088 -1381 -1057
rect 1381 -1088 1398 -1057
rect -1398 -1105 -1350 -1088
rect 1350 -1105 1398 -1088
<< viali >>
rect -1350 1088 1350 1105
rect -1398 -1057 -1381 1057
rect -1300 1019 -816 1036
rect -771 1019 -287 1036
rect -242 1019 242 1036
rect 287 1019 771 1036
rect 816 1019 1300 1036
rect -1331 -994 -1314 994
rect -802 -994 -785 994
rect -273 -994 -256 994
rect 256 -994 273 994
rect 785 -994 802 994
rect 1314 -994 1331 994
rect -1300 -1036 -816 -1019
rect -771 -1036 -287 -1019
rect -242 -1036 242 -1019
rect 287 -1036 771 -1019
rect 816 -1036 1300 -1019
rect 1381 -1057 1398 1057
rect -1350 -1105 1350 -1088
<< metal1 >>
rect -1404 1105 1404 1111
rect -1404 1088 -1350 1105
rect 1350 1088 1404 1105
rect -1404 1082 1404 1088
rect -1404 1057 -1375 1082
rect -1404 -1057 -1398 1057
rect -1381 950 -1375 1057
rect 1375 1057 1404 1082
rect -1308 1045 1308 1048
rect -1308 1019 -1305 1045
rect 1305 1019 1308 1045
rect -1308 1016 1308 1019
rect -1334 994 -1311 1000
rect -1334 950 -1331 994
rect -1381 850 -1331 950
rect -1381 750 -1375 850
rect -1334 750 -1331 850
rect -1381 650 -1331 750
rect -1381 550 -1375 650
rect -1334 550 -1331 650
rect -1381 450 -1331 550
rect -1381 350 -1375 450
rect -1334 350 -1331 450
rect -1381 250 -1331 350
rect -1381 150 -1375 250
rect -1334 150 -1331 250
rect -1381 50 -1331 150
rect -1381 -50 -1375 50
rect -1334 -50 -1331 50
rect -1381 -150 -1331 -50
rect -1381 -250 -1375 -150
rect -1334 -250 -1331 -150
rect -1381 -350 -1331 -250
rect -1381 -450 -1375 -350
rect -1334 -450 -1331 -350
rect -1381 -550 -1331 -450
rect -1381 -650 -1375 -550
rect -1334 -650 -1331 -550
rect -1381 -750 -1331 -650
rect -1381 -850 -1375 -750
rect -1334 -850 -1331 -750
rect -1381 -950 -1331 -850
rect -1381 -1057 -1375 -950
rect -1334 -994 -1331 -950
rect -1314 950 -1311 994
rect -805 994 -782 1000
rect -805 950 -802 994
rect -1314 850 -802 950
rect -1314 750 -1311 850
rect -805 750 -802 850
rect -1314 650 -802 750
rect -1314 550 -1311 650
rect -805 550 -802 650
rect -1314 450 -802 550
rect -1314 350 -1311 450
rect -805 350 -802 450
rect -1314 250 -802 350
rect -1314 150 -1311 250
rect -805 150 -802 250
rect -1314 50 -802 150
rect -1314 -50 -1311 50
rect -805 -50 -802 50
rect -1314 -150 -802 -50
rect -1314 -250 -1311 -150
rect -805 -250 -802 -150
rect -1314 -350 -802 -250
rect -1314 -450 -1311 -350
rect -805 -450 -802 -350
rect -1314 -550 -802 -450
rect -1314 -650 -1311 -550
rect -805 -650 -802 -550
rect -1314 -750 -802 -650
rect -1314 -850 -1311 -750
rect -805 -850 -802 -750
rect -1314 -950 -802 -850
rect -1314 -994 -1311 -950
rect -1334 -1000 -1311 -994
rect -805 -994 -802 -950
rect -785 950 -782 994
rect -276 994 -253 1000
rect -276 950 -273 994
rect -785 850 -273 950
rect -785 750 -782 850
rect -276 750 -273 850
rect -785 650 -273 750
rect -785 550 -782 650
rect -276 550 -273 650
rect -785 450 -273 550
rect -785 350 -782 450
rect -276 350 -273 450
rect -785 250 -273 350
rect -785 150 -782 250
rect -276 150 -273 250
rect -785 50 -273 150
rect -785 -50 -782 50
rect -276 -50 -273 50
rect -785 -150 -273 -50
rect -785 -250 -782 -150
rect -276 -250 -273 -150
rect -785 -350 -273 -250
rect -785 -450 -782 -350
rect -276 -450 -273 -350
rect -785 -550 -273 -450
rect -785 -650 -782 -550
rect -276 -650 -273 -550
rect -785 -750 -273 -650
rect -785 -850 -782 -750
rect -276 -850 -273 -750
rect -785 -950 -273 -850
rect -785 -994 -782 -950
rect -805 -1000 -782 -994
rect -276 -994 -273 -950
rect -256 950 -253 994
rect 253 994 276 1000
rect 253 950 256 994
rect -256 850 256 950
rect -256 750 -253 850
rect 253 750 256 850
rect -256 650 256 750
rect -256 550 -253 650
rect 253 550 256 650
rect -256 450 256 550
rect -256 350 -253 450
rect 253 350 256 450
rect -256 250 256 350
rect -256 150 -253 250
rect 253 150 256 250
rect -256 50 256 150
rect -256 -50 -253 50
rect 253 -50 256 50
rect -256 -150 256 -50
rect -256 -250 -253 -150
rect 253 -250 256 -150
rect -256 -350 256 -250
rect -256 -450 -253 -350
rect 253 -450 256 -350
rect -256 -550 256 -450
rect -256 -650 -253 -550
rect 253 -650 256 -550
rect -256 -750 256 -650
rect -256 -850 -253 -750
rect 253 -850 256 -750
rect -256 -950 256 -850
rect -256 -994 -253 -950
rect -276 -1000 -253 -994
rect 253 -994 256 -950
rect 273 950 276 994
rect 782 994 805 1000
rect 782 950 785 994
rect 273 850 785 950
rect 273 750 276 850
rect 782 750 785 850
rect 273 650 785 750
rect 273 550 276 650
rect 782 550 785 650
rect 273 450 785 550
rect 273 350 276 450
rect 782 350 785 450
rect 273 250 785 350
rect 273 150 276 250
rect 782 150 785 250
rect 273 50 785 150
rect 273 -50 276 50
rect 782 -50 785 50
rect 273 -150 785 -50
rect 273 -250 276 -150
rect 782 -250 785 -150
rect 273 -350 785 -250
rect 273 -450 276 -350
rect 782 -450 785 -350
rect 273 -550 785 -450
rect 273 -650 276 -550
rect 782 -650 785 -550
rect 273 -750 785 -650
rect 273 -850 276 -750
rect 782 -850 785 -750
rect 273 -950 785 -850
rect 273 -994 276 -950
rect 253 -1000 276 -994
rect 782 -994 785 -950
rect 802 950 805 994
rect 1311 994 1334 1000
rect 1311 950 1314 994
rect 802 850 1314 950
rect 802 750 805 850
rect 1311 750 1314 850
rect 802 650 1314 750
rect 802 550 805 650
rect 1311 550 1314 650
rect 802 450 1314 550
rect 802 350 805 450
rect 1311 350 1314 450
rect 802 250 1314 350
rect 802 150 805 250
rect 1311 150 1314 250
rect 802 50 1314 150
rect 802 -50 805 50
rect 1311 -50 1314 50
rect 802 -150 1314 -50
rect 802 -250 805 -150
rect 1311 -250 1314 -150
rect 802 -350 1314 -250
rect 802 -450 805 -350
rect 1311 -450 1314 -350
rect 802 -550 1314 -450
rect 802 -650 805 -550
rect 1311 -650 1314 -550
rect 802 -750 1314 -650
rect 802 -850 805 -750
rect 1311 -850 1314 -750
rect 802 -950 1314 -850
rect 802 -994 805 -950
rect 782 -1000 805 -994
rect 1311 -994 1314 -950
rect 1331 950 1334 994
rect 1375 950 1381 1057
rect 1331 850 1381 950
rect 1331 750 1334 850
rect 1375 750 1381 850
rect 1331 650 1381 750
rect 1331 550 1334 650
rect 1375 550 1381 650
rect 1331 450 1381 550
rect 1331 350 1334 450
rect 1375 350 1381 450
rect 1331 250 1381 350
rect 1331 150 1334 250
rect 1375 150 1381 250
rect 1331 50 1381 150
rect 1331 -50 1334 50
rect 1375 -50 1381 50
rect 1331 -150 1381 -50
rect 1331 -250 1334 -150
rect 1375 -250 1381 -150
rect 1331 -350 1381 -250
rect 1331 -450 1334 -350
rect 1375 -450 1381 -350
rect 1331 -550 1381 -450
rect 1331 -650 1334 -550
rect 1375 -650 1381 -550
rect 1331 -750 1381 -650
rect 1331 -850 1334 -750
rect 1375 -850 1381 -750
rect 1331 -950 1381 -850
rect 1331 -994 1334 -950
rect 1311 -1000 1334 -994
rect -1308 -1019 1308 -1016
rect -1308 -1045 -1305 -1019
rect 1305 -1045 1308 -1019
rect -1308 -1048 1308 -1045
rect -1404 -1082 -1375 -1057
rect 1375 -1057 1381 -950
rect 1398 -1057 1404 1057
rect 1375 -1082 1404 -1057
rect -1404 -1088 1404 -1082
rect -1404 -1105 -1350 -1088
rect 1350 -1105 1404 -1088
rect -1404 -1111 1404 -1105
<< via1 >>
rect -1305 1036 1305 1045
rect -1305 1019 -1300 1036
rect -1300 1019 -816 1036
rect -816 1019 -771 1036
rect -771 1019 -287 1036
rect -287 1019 -242 1036
rect -242 1019 242 1036
rect 242 1019 287 1036
rect 287 1019 771 1036
rect 771 1019 816 1036
rect 816 1019 1300 1036
rect 1300 1019 1305 1036
rect -1305 -1036 -1300 -1019
rect -1300 -1036 -816 -1019
rect -816 -1036 -771 -1019
rect -771 -1036 -287 -1019
rect -287 -1036 -242 -1019
rect -242 -1036 242 -1019
rect 242 -1036 287 -1019
rect 287 -1036 771 -1019
rect 771 -1036 816 -1019
rect 816 -1036 1300 -1019
rect 1300 -1036 1305 -1019
rect -1305 -1045 1305 -1036
<< metal2 >>
rect -1308 1045 1308 1066
rect -1308 1019 -1305 1045
rect 1305 1019 1308 1045
rect -1308 1016 1308 1019
rect -1308 -1019 1308 -1016
rect -1308 -1045 -1305 -1019
rect 1305 -1045 1308 -1019
rect -1308 -1066 1308 -1045
<< properties >>
string FIXED_BBOX -1389 -1096 1389 1096
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 20 l 5 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
