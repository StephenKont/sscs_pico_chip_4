magic
tech sky130A
magscale 1 2
timestamp 1667842615
<< viali >>
rect 3186 7076 3220 7110
rect 3328 7076 3362 7110
rect 3408 7076 3442 7110
rect 3494 7076 3528 7110
rect 3578 7076 3612 7110
rect 3650 7076 3684 7110
rect 6384 7078 6418 7112
rect 6566 7076 6600 7110
rect 6698 7076 6732 7110
rect 6960 7076 6994 7110
rect 7086 7076 7120 7110
rect 7180 7076 7214 7110
rect 4134 1992 4170 2028
rect 4232 1994 4268 2030
rect 4344 1994 4380 2030
rect 4430 1992 4466 2028
<< metal1 >>
rect 6122 8148 6240 8152
rect 3722 8080 6240 8148
rect 758 7720 1036 7760
rect 758 7566 812 7720
rect 984 7566 1036 7720
rect 758 7238 1036 7566
rect 3724 7270 3800 8080
rect 6122 7814 6240 8080
rect 6076 7770 6280 7814
rect 6076 7718 6102 7770
rect 6256 7718 6280 7770
rect 6076 7702 6280 7718
rect 10624 7328 14546 7378
rect 3524 7216 4060 7270
rect 6950 7268 7226 7276
rect 10624 7268 10684 7328
rect 6950 7218 10684 7268
rect 6950 7158 7226 7218
rect 3176 7112 7228 7158
rect 3176 7110 6384 7112
rect 3176 7076 3186 7110
rect 3220 7076 3328 7110
rect 3362 7076 3408 7110
rect 3442 7076 3494 7110
rect 3528 7076 3578 7110
rect 3612 7076 3650 7110
rect 3684 7078 6384 7110
rect 6418 7110 7228 7112
rect 6418 7078 6566 7110
rect 3684 7076 6566 7078
rect 6600 7076 6698 7110
rect 6732 7076 6960 7110
rect 6994 7076 7086 7110
rect 7120 7076 7180 7110
rect 7214 7076 7228 7110
rect 3176 7042 7228 7076
rect 6950 7040 7004 7042
rect 7078 7040 7128 7042
rect 7168 7040 7226 7042
rect 184 6000 252 6008
rect 184 5994 192 6000
rect -508 5952 192 5994
rect 184 5948 192 5952
rect 244 5948 252 6000
rect 184 5942 252 5948
rect 14496 5266 14546 7328
rect 11146 5216 14546 5266
rect 14014 3972 14084 4030
rect 14014 3920 14022 3972
rect 14074 3920 14084 3972
rect 14014 3896 14084 3920
rect 4150 2198 4502 2210
rect 4150 2194 4310 2198
rect 4468 2194 4502 2198
rect 408 2184 1868 2194
rect 408 2132 414 2184
rect 466 2132 1868 2184
rect 408 2124 1868 2132
rect 4150 2122 4160 2194
rect 4486 2122 4502 2194
rect 4150 2114 4502 2122
rect 4108 2036 4488 2074
rect 10074 2036 10124 3100
rect 14496 3098 14546 5216
rect 10620 3048 14546 3098
rect 4108 2030 10124 2036
rect 4108 2028 4232 2030
rect 4108 1992 4134 2028
rect 4170 1994 4232 2028
rect 4268 1994 4344 2030
rect 4380 2028 10124 2030
rect 4380 1994 4430 2028
rect 4170 1992 4430 1994
rect 4466 1992 10124 2028
rect 4108 1986 10124 1992
rect 4108 1956 4488 1986
rect 4122 1954 4488 1956
<< via1 >>
rect 812 7566 984 7720
rect 6102 7718 6256 7770
rect 14024 6902 14076 6954
rect 192 5948 244 6000
rect 14022 3920 14074 3972
rect 4310 2194 4468 2198
rect 414 2132 466 2184
rect 4160 2122 4486 2194
<< metal2 >>
rect 14012 8524 14084 8530
rect -1918 8452 14084 8524
rect -1916 7402 -354 8452
rect 6076 7770 6280 7814
rect 788 7732 1006 7744
rect 266 7660 726 7662
rect 788 7660 800 7732
rect 88 7598 800 7660
rect 88 -4668 152 7598
rect 186 7596 800 7598
rect 788 7554 800 7596
rect 994 7554 1006 7732
rect 6076 7718 6102 7770
rect 6256 7718 6280 7770
rect 6076 7702 6280 7718
rect 788 7542 1006 7554
rect 14012 6988 14084 8452
rect 14014 6954 14084 6988
rect 14014 6902 14024 6954
rect 14076 6902 14084 6954
rect 184 6000 252 6008
rect 184 5948 192 6000
rect 244 5948 252 6000
rect 184 5942 252 5948
rect 414 2194 464 5966
rect 14014 3972 14084 6902
rect 14014 3920 14022 3972
rect 14074 3920 14084 3972
rect 14014 3896 14084 3920
rect 4230 2212 4512 2236
rect 4230 2210 4242 2212
rect 4150 2194 4242 2210
rect 408 2184 470 2194
rect 408 2132 414 2184
rect 466 2132 470 2184
rect 408 2124 470 2132
rect 4150 2122 4160 2194
rect 4496 2142 4512 2212
rect 4486 2126 4512 2142
rect 4486 2122 4502 2126
rect 4150 2114 4502 2122
rect -8946 -5358 636 -5306
rect -8946 -5704 -34 -5358
rect 196 -5704 636 -5358
rect -8946 -6020 -32 -5704
rect 188 -6020 636 -5704
rect -8946 -7010 636 -6020
<< via2 >>
rect 800 7720 994 7732
rect 800 7566 812 7720
rect 812 7566 984 7720
rect 984 7566 994 7720
rect 800 7554 994 7566
rect 4242 2198 4496 2212
rect 4242 2194 4310 2198
rect 4310 2194 4468 2198
rect 4468 2194 4496 2198
rect 4242 2142 4486 2194
rect 4486 2142 4496 2194
rect 4306 2136 4474 2142
rect -34 -5704 196 -5358
rect -32 -6020 188 -5704
<< metal3 >>
rect 776 7732 1036 7746
rect 776 7554 800 7732
rect 994 7554 1036 7732
rect 776 7536 1036 7554
rect 776 7534 952 7536
rect 4180 2360 4620 2378
rect 4180 2126 4196 2360
rect 4608 2126 4620 2360
rect 4180 2116 4620 2126
rect -238 -5330 722 -5308
rect -240 -5358 1306 -5330
rect -240 -5496 -34 -5358
rect -240 -6784 -120 -5496
rect 196 -5704 1306 -5358
rect 188 -6020 1306 -5704
rect 166 -6784 1306 -6020
rect -240 -6816 1306 -6784
rect -242 -6962 1306 -6816
rect -242 -7010 688 -6962
<< via3 >>
rect 4196 2212 4608 2360
rect 4196 2142 4242 2212
rect 4242 2142 4496 2212
rect 4496 2142 4608 2212
rect 4196 2136 4306 2142
rect 4306 2136 4474 2142
rect 4474 2136 4608 2142
rect 4196 2126 4608 2136
rect -120 -5704 -34 -5496
rect -34 -5704 166 -5496
rect -120 -6020 -32 -5704
rect -32 -6020 166 -5704
rect -120 -6784 166 -6020
<< metal4 >>
rect 4160 2360 4642 2380
rect 4160 2126 4196 2360
rect 4608 2126 4642 2360
rect 4160 1658 4642 2126
<< via4 >>
rect -156 -5496 242 -5458
rect -156 -6784 -120 -5496
rect -120 -6784 166 -5496
rect 166 -6784 242 -5496
rect -156 -6830 242 -6784
<< metal5 >>
rect -156 -5362 244 -5334
rect -220 -5366 244 -5362
rect -220 -5458 872 -5366
rect -220 -6830 -156 -5458
rect 242 -6830 872 -5458
rect -220 -6880 872 -6830
rect -130 -6882 872 -6880
use current_source  current_source_0
timestamp 1667842615
transform 1 0 3796 0 1 1152
box -1962 1810 10276 3598
use op_amp_layout1  op_amp_layout1_0
timestamp 1666558548
transform 1 0 4626 0 1 1602
box -4388 1254 9738 6166
use pass_element  pass_element_0
timestamp 1666808413
transform 0 1 -20554 -1 0 9064
box 1242 11596 14806 20746
use sky130_fd_pr__cap_mim_m3_1_3VRXMH  sky130_fd_pr__cap_mim_m3_1_3VRXMH_0
timestamp 1666550119
transform 0 -1 7870 1 0 -3773
box -4909 -7450 5525 7456
use sky130_fd_pr__res_high_po_0p35_8W29VJ  sky130_fd_pr__res_high_po_0p35_8W29VJ_0
timestamp 1666532281
transform 0 -1 2145 1 0 7241
box -201 -1571 201 1571
use sky130_fd_pr__res_high_po_0p35_8W29VJ  sky130_fd_pr__res_high_po_0p35_8W29VJ_1
timestamp 1666532281
transform 0 -1 3083 1 0 2159
box -201 -1571 201 1571
use sky130_fd_pr__res_high_po_0p35_V8E24B  sky130_fd_pr__res_high_po_0p35_V8E24B_0
timestamp 1666532426
transform 0 1 5648 -1 0 7241
box -201 -1812 201 1812
<< labels >>
rlabel metal1 812 7364 984 7518 1 Vout
rlabel metal2 -1728 7962 -568 8416 1 VDD
rlabel space 9750 7710 9922 7760 1 Vref
<< end >>
