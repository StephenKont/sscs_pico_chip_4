magic
tech sky130A
magscale 1 2
timestamp 1666553439
<< metal3 >>
rect -18947 3444 -12709 6250
rect -12488 3444 -6253 6250
rect -5889 3444 349 6250
rect 850 3444 7089 6250
rect 7449 3444 13687 6250
rect 14048 3444 20347 6250
rect -18947 2844 20347 3444
rect -18947 50 -12709 2844
rect -12488 2818 349 2844
rect -12488 50 -6253 2818
rect -5889 50 349 2818
rect 850 50 7089 2844
rect 7449 50 13687 2844
rect 14048 50 20347 2844
rect -15909 -50 -15775 50
rect -9451 -50 -9317 50
rect -2853 -50 -2719 50
rect 3883 -50 4017 50
rect 10483 -50 10617 50
rect 17083 -50 17217 50
rect -18947 -2806 -12709 -50
rect -12488 -2806 -6253 -50
rect -5889 -2806 349 -50
rect 850 -2806 7089 -50
rect 7449 -2806 13687 -50
rect 14048 -2806 20347 -50
rect -18947 -3406 20347 -2806
rect -18947 -6250 -12709 -3406
rect -12488 -3414 20347 -3406
rect -12488 -6250 -6253 -3414
rect -5889 -3418 20347 -3414
rect -5889 -6250 349 -3418
rect 850 -3442 20347 -3418
rect 850 -3534 13687 -3442
rect 850 -6250 7089 -3534
rect 7449 -6250 13687 -3534
rect 14048 -6250 20347 -3442
<< mimcap >>
rect -18847 6110 -12847 6150
rect -18847 190 -18807 6110
rect -12887 190 -12847 6110
rect -18847 150 -12847 190
rect -12388 6110 -6388 6150
rect -12388 190 -12348 6110
rect -6428 190 -6388 6110
rect -12388 150 -6388 190
rect -5789 6110 211 6150
rect -5789 190 -5749 6110
rect 171 190 211 6110
rect -5789 150 211 190
rect 950 6110 6950 6150
rect 950 190 990 6110
rect 6910 190 6950 6110
rect 950 150 6950 190
rect 7549 6110 13549 6150
rect 7549 190 7589 6110
rect 13509 190 13549 6110
rect 7549 150 13549 190
rect 14148 6110 20148 6150
rect 14148 190 14188 6110
rect 20108 190 20148 6110
rect 14148 150 20148 190
rect -18847 -190 -12847 -150
rect -18847 -6110 -18807 -190
rect -12887 -6110 -12847 -190
rect -18847 -6150 -12847 -6110
rect -12388 -190 -6388 -150
rect -12388 -6110 -12348 -190
rect -6428 -6110 -6388 -190
rect -12388 -6150 -6388 -6110
rect -5789 -190 211 -150
rect -5789 -6110 -5749 -190
rect 171 -6110 211 -190
rect -5789 -6150 211 -6110
rect 950 -190 6950 -150
rect 950 -6110 990 -190
rect 6910 -6110 6950 -190
rect 950 -6150 6950 -6110
rect 7549 -190 13549 -150
rect 7549 -6110 7589 -190
rect 13509 -6110 13549 -190
rect 7549 -6150 13549 -6110
rect 14148 -190 20148 -150
rect 14148 -6110 14188 -190
rect 20108 -6110 20148 -190
rect 14148 -6150 20148 -6110
<< mimcapcontact >>
rect -18807 190 -12887 6110
rect -12348 190 -6428 6110
rect -5749 190 171 6110
rect 990 190 6910 6110
rect 7589 190 13509 6110
rect 14188 190 20108 6110
rect -18807 -6110 -12887 -190
rect -12348 -6110 -6428 -190
rect -5749 -6110 171 -190
rect 990 -6110 6910 -190
rect 7589 -6110 13509 -190
rect 14188 -6110 20108 -190
<< metal4 >>
rect -15899 6111 -15795 6300
rect -9440 6111 -9336 6300
rect -2841 6111 -2737 6300
rect 3898 6111 4002 6300
rect 10497 6111 10601 6300
rect 17096 6111 17200 6300
rect -18808 6110 -12886 6111
rect -18808 190 -18807 6110
rect -12887 3444 -12886 6110
rect -12349 6110 -6427 6111
rect -12349 3444 -12348 6110
rect -12887 2844 -12348 3444
rect -12887 190 -12886 2844
rect -18808 189 -12886 190
rect -12349 190 -12348 2844
rect -6428 3444 -6427 6110
rect -5750 6110 172 6111
rect -5750 3444 -5749 6110
rect -6428 2818 -5749 3444
rect -6428 190 -6427 2818
rect -12349 189 -6427 190
rect -5750 190 -5749 2818
rect 171 3444 172 6110
rect 989 6110 6911 6111
rect 989 3444 990 6110
rect 171 2844 990 3444
rect 171 190 172 2844
rect -5750 189 172 190
rect 989 190 990 2844
rect 6910 3444 6911 6110
rect 7588 6110 13510 6111
rect 7588 3444 7589 6110
rect 6910 2844 7589 3444
rect 6910 190 6911 2844
rect 989 189 6911 190
rect 7588 190 7589 2844
rect 13509 3444 13510 6110
rect 14187 6110 20109 6111
rect 14187 3444 14188 6110
rect 13509 2844 14188 3444
rect 13509 190 13510 2844
rect 7588 189 13510 190
rect 14187 190 14188 2844
rect 20108 190 20109 6110
rect 14187 189 20109 190
rect -15899 -189 -15795 189
rect -9440 -189 -9336 189
rect -2841 -189 -2737 189
rect 3898 -189 4002 189
rect 10497 -189 10601 189
rect 17096 -189 17200 189
rect -18808 -190 -12886 -189
rect -18808 -6110 -18807 -190
rect -12887 -2806 -12886 -190
rect -12349 -190 -6427 -189
rect -12349 -2806 -12348 -190
rect -12887 -3406 -12348 -2806
rect -12887 -6110 -12886 -3406
rect -18808 -6111 -12886 -6110
rect -12349 -6110 -12348 -3406
rect -6428 -2806 -6427 -190
rect -5750 -190 172 -189
rect -5750 -2806 -5749 -190
rect -6428 -3414 -5749 -2806
rect -6428 -6110 -6427 -3414
rect -12349 -6111 -6427 -6110
rect -5750 -6110 -5749 -3414
rect 171 -2806 172 -190
rect 989 -190 6911 -189
rect 989 -2806 990 -190
rect 171 -3418 990 -2806
rect 171 -6110 172 -3418
rect -5750 -6111 172 -6110
rect 989 -6110 990 -3418
rect 6910 -2806 6911 -190
rect 7588 -190 13510 -189
rect 7588 -2806 7589 -190
rect 6910 -3534 7589 -2806
rect 6910 -6110 6911 -3534
rect 989 -6111 6911 -6110
rect 7588 -6110 7589 -3534
rect 13509 -2806 13510 -190
rect 14187 -190 20109 -189
rect 14187 -2806 14188 -190
rect 13509 -3442 14188 -2806
rect 13509 -6110 13510 -3442
rect 7588 -6111 13510 -6110
rect 14187 -6110 14188 -3442
rect 20108 -6110 20109 -190
rect 14187 -6111 20109 -6110
rect -15899 -6300 -15795 -6111
rect -9440 -6300 -9336 -6111
rect -2841 -6300 -2737 -6111
rect 3898 -6300 4002 -6111
rect 10497 -6300 10601 -6111
rect 17096 -6300 17200 -6111
<< properties >>
string FIXED_BBOX 12648 50 18848 6250
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 6 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
