magic
tech sky130A
magscale 1 2
timestamp 1666554250
<< nwell >>
rect -807 -719 807 719
<< pmoslvt >>
rect -611 -500 -541 500
rect -483 -500 -413 500
rect -355 -500 -285 500
rect -227 -500 -157 500
rect -99 -500 -29 500
rect 29 -500 99 500
rect 157 -500 227 500
rect 285 -500 355 500
rect 413 -500 483 500
rect 541 -500 611 500
<< pdiff >>
rect -669 488 -611 500
rect -669 -488 -657 488
rect -623 -488 -611 488
rect -669 -500 -611 -488
rect -541 488 -483 500
rect -541 -488 -529 488
rect -495 -488 -483 488
rect -541 -500 -483 -488
rect -413 488 -355 500
rect -413 -488 -401 488
rect -367 -488 -355 488
rect -413 -500 -355 -488
rect -285 488 -227 500
rect -285 -488 -273 488
rect -239 -488 -227 488
rect -285 -500 -227 -488
rect -157 488 -99 500
rect -157 -488 -145 488
rect -111 -488 -99 488
rect -157 -500 -99 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 99 488 157 500
rect 99 -488 111 488
rect 145 -488 157 488
rect 99 -500 157 -488
rect 227 488 285 500
rect 227 -488 239 488
rect 273 -488 285 488
rect 227 -500 285 -488
rect 355 488 413 500
rect 355 -488 367 488
rect 401 -488 413 488
rect 355 -500 413 -488
rect 483 488 541 500
rect 483 -488 495 488
rect 529 -488 541 488
rect 483 -500 541 -488
rect 611 488 669 500
rect 611 -488 623 488
rect 657 -488 669 488
rect 611 -500 669 -488
<< pdiffc >>
rect -657 -488 -623 488
rect -529 -488 -495 488
rect -401 -488 -367 488
rect -273 -488 -239 488
rect -145 -488 -111 488
rect -17 -488 17 488
rect 111 -488 145 488
rect 239 -488 273 488
rect 367 -488 401 488
rect 495 -488 529 488
rect 623 -488 657 488
<< nsubdiff >>
rect -771 649 -675 683
rect 675 649 771 683
rect -771 587 -737 649
rect 737 587 771 649
rect -771 -649 -737 -587
rect 737 -649 771 -587
rect -771 -683 -675 -649
rect 675 -683 771 -649
<< nsubdiffcont >>
rect -675 649 675 683
rect -771 -587 -737 587
rect 737 -587 771 587
rect -675 -683 675 -649
<< poly >>
rect -611 581 -541 597
rect -611 547 -595 581
rect -557 547 -541 581
rect -611 500 -541 547
rect -483 581 -413 597
rect -483 547 -467 581
rect -429 547 -413 581
rect -483 500 -413 547
rect -355 581 -285 597
rect -355 547 -339 581
rect -301 547 -285 581
rect -355 500 -285 547
rect -227 581 -157 597
rect -227 547 -211 581
rect -173 547 -157 581
rect -227 500 -157 547
rect -99 581 -29 597
rect -99 547 -83 581
rect -45 547 -29 581
rect -99 500 -29 547
rect 29 581 99 597
rect 29 547 45 581
rect 83 547 99 581
rect 29 500 99 547
rect 157 581 227 597
rect 157 547 173 581
rect 211 547 227 581
rect 157 500 227 547
rect 285 581 355 597
rect 285 547 301 581
rect 339 547 355 581
rect 285 500 355 547
rect 413 581 483 597
rect 413 547 429 581
rect 467 547 483 581
rect 413 500 483 547
rect 541 581 611 597
rect 541 547 557 581
rect 595 547 611 581
rect 541 500 611 547
rect -611 -547 -541 -500
rect -611 -581 -595 -547
rect -557 -581 -541 -547
rect -611 -597 -541 -581
rect -483 -547 -413 -500
rect -483 -581 -467 -547
rect -429 -581 -413 -547
rect -483 -597 -413 -581
rect -355 -547 -285 -500
rect -355 -581 -339 -547
rect -301 -581 -285 -547
rect -355 -597 -285 -581
rect -227 -547 -157 -500
rect -227 -581 -211 -547
rect -173 -581 -157 -547
rect -227 -597 -157 -581
rect -99 -547 -29 -500
rect -99 -581 -83 -547
rect -45 -581 -29 -547
rect -99 -597 -29 -581
rect 29 -547 99 -500
rect 29 -581 45 -547
rect 83 -581 99 -547
rect 29 -597 99 -581
rect 157 -547 227 -500
rect 157 -581 173 -547
rect 211 -581 227 -547
rect 157 -597 227 -581
rect 285 -547 355 -500
rect 285 -581 301 -547
rect 339 -581 355 -547
rect 285 -597 355 -581
rect 413 -547 483 -500
rect 413 -581 429 -547
rect 467 -581 483 -547
rect 413 -597 483 -581
rect 541 -547 611 -500
rect 541 -581 557 -547
rect 595 -581 611 -547
rect 541 -597 611 -581
<< polycont >>
rect -595 547 -557 581
rect -467 547 -429 581
rect -339 547 -301 581
rect -211 547 -173 581
rect -83 547 -45 581
rect 45 547 83 581
rect 173 547 211 581
rect 301 547 339 581
rect 429 547 467 581
rect 557 547 595 581
rect -595 -581 -557 -547
rect -467 -581 -429 -547
rect -339 -581 -301 -547
rect -211 -581 -173 -547
rect -83 -581 -45 -547
rect 45 -581 83 -547
rect 173 -581 211 -547
rect 301 -581 339 -547
rect 429 -581 467 -547
rect 557 -581 595 -547
<< locali >>
rect -771 649 -675 683
rect 675 649 771 683
rect -771 587 -737 649
rect 737 587 771 649
rect -611 547 -595 581
rect -557 547 -541 581
rect -483 547 -467 581
rect -429 547 -413 581
rect -355 547 -339 581
rect -301 547 -285 581
rect -227 547 -211 581
rect -173 547 -157 581
rect -99 547 -83 581
rect -45 547 -29 581
rect 29 547 45 581
rect 83 547 99 581
rect 157 547 173 581
rect 211 547 227 581
rect 285 547 301 581
rect 339 547 355 581
rect 413 547 429 581
rect 467 547 483 581
rect 541 547 557 581
rect 595 547 611 581
rect -657 488 -623 504
rect -657 -504 -623 -488
rect -529 488 -495 504
rect -529 -504 -495 -488
rect -401 488 -367 504
rect -401 -504 -367 -488
rect -273 488 -239 504
rect -273 -504 -239 -488
rect -145 488 -111 504
rect -145 -504 -111 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 111 488 145 504
rect 111 -504 145 -488
rect 239 488 273 504
rect 239 -504 273 -488
rect 367 488 401 504
rect 367 -504 401 -488
rect 495 488 529 504
rect 495 -504 529 -488
rect 623 488 657 504
rect 623 -504 657 -488
rect -611 -581 -595 -547
rect -557 -581 -541 -547
rect -483 -581 -467 -547
rect -429 -581 -413 -547
rect -355 -581 -339 -547
rect -301 -581 -285 -547
rect -227 -581 -211 -547
rect -173 -581 -157 -547
rect -99 -581 -83 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 83 -581 99 -547
rect 157 -581 173 -547
rect 211 -581 227 -547
rect 285 -581 301 -547
rect 339 -581 355 -547
rect 413 -581 429 -547
rect 467 -581 483 -547
rect 541 -581 557 -547
rect 595 -581 611 -547
rect -771 -649 -737 -587
rect 737 -649 771 -587
rect -771 -683 -675 -649
rect 675 -683 771 -649
<< viali >>
rect -595 547 -557 581
rect -467 547 -429 581
rect -339 547 -301 581
rect -211 547 -173 581
rect -83 547 -45 581
rect 45 547 83 581
rect 173 547 211 581
rect 301 547 339 581
rect 429 547 467 581
rect 557 547 595 581
rect -657 -488 -623 488
rect -529 -488 -495 488
rect -401 -488 -367 488
rect -273 -488 -239 488
rect -145 -488 -111 488
rect -17 -488 17 488
rect 111 -488 145 488
rect 239 -488 273 488
rect 367 -488 401 488
rect 495 -488 529 488
rect 623 -488 657 488
rect -595 -581 -557 -547
rect -467 -581 -429 -547
rect -339 -581 -301 -547
rect -211 -581 -173 -547
rect -83 -581 -45 -547
rect 45 -581 83 -547
rect 173 -581 211 -547
rect 301 -581 339 -547
rect 429 -581 467 -547
rect 557 -581 595 -547
<< metal1 >>
rect -611 581 611 597
rect -611 547 -595 581
rect -557 547 -467 581
rect -429 547 -339 581
rect -301 547 -211 581
rect -173 547 -83 581
rect -45 547 45 581
rect 83 547 173 581
rect 211 547 301 581
rect 339 547 429 581
rect 467 547 557 581
rect 595 547 611 581
rect -611 541 611 547
rect -663 488 -617 500
rect -663 -488 -657 488
rect -623 -488 -617 488
rect -663 -500 -617 -488
rect -535 488 -489 500
rect -535 -488 -529 488
rect -495 -488 -489 488
rect -535 -500 -489 -488
rect -407 488 -361 500
rect -407 -488 -401 488
rect -367 -488 -361 488
rect -407 -500 -361 -488
rect -279 488 -233 500
rect -279 -488 -273 488
rect -239 -488 -233 488
rect -279 -500 -233 -488
rect -151 488 -105 500
rect -151 -488 -145 488
rect -111 -488 -105 488
rect -151 -500 -105 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 105 488 151 500
rect 105 -488 111 488
rect 145 -488 151 488
rect 105 -500 151 -488
rect 233 488 279 500
rect 233 -488 239 488
rect 273 -488 279 488
rect 233 -500 279 -488
rect 361 488 407 500
rect 361 -488 367 488
rect 401 -488 407 488
rect 361 -500 407 -488
rect 489 488 535 500
rect 489 -488 495 488
rect 529 -488 535 488
rect 489 -500 535 -488
rect 617 488 663 500
rect 617 -488 623 488
rect 657 -488 663 488
rect 617 -500 663 -488
rect -611 -547 611 -541
rect -611 -581 -595 -547
rect -557 -581 -467 -547
rect -429 -581 -339 -547
rect -301 -581 -211 -547
rect -173 -581 -83 -547
rect -45 -581 45 -547
rect 83 -581 173 -547
rect 211 -581 301 -547
rect 339 -581 429 -547
rect 467 -581 557 -547
rect 595 -581 611 -547
rect -611 -597 611 -581
<< properties >>
string FIXED_BBOX -754 -666 754 666
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5 l 0.35 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
