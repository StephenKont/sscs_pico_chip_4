magic
tech sky130A
magscale 1 2
timestamp 1668293870
<< nwell >>
rect -321 -319 321 319
<< pmos >>
rect -125 -100 125 100
<< pdiff >>
rect -183 88 -125 100
rect -183 -88 -171 88
rect -137 -88 -125 88
rect -183 -100 -125 -88
rect 125 88 183 100
rect 125 -88 137 88
rect 171 -88 183 88
rect 125 -100 183 -88
<< pdiffc >>
rect -171 -88 -137 88
rect 137 -88 171 88
<< nsubdiff >>
rect -285 249 -189 283
rect 189 249 285 283
rect -285 187 -251 249
rect 251 187 285 249
rect -285 -249 -251 -187
rect 251 -249 285 -187
rect -285 -283 -189 -249
rect 189 -283 285 -249
<< nsubdiffcont >>
rect -189 249 189 283
rect -285 -187 -251 187
rect 251 -187 285 187
rect -189 -283 189 -249
<< poly >>
rect -125 181 125 197
rect -125 147 -109 181
rect 109 147 125 181
rect -125 100 125 147
rect -125 -147 125 -100
rect -125 -181 -109 -147
rect 109 -181 125 -147
rect -125 -197 125 -181
<< polycont >>
rect -109 147 109 181
rect -109 -181 109 -147
<< locali >>
rect -285 249 -189 283
rect 189 249 285 283
rect -285 187 -251 249
rect 251 187 285 249
rect -125 147 -109 181
rect 109 147 125 181
rect -171 88 -137 104
rect -171 -104 -137 -88
rect 137 88 171 104
rect 137 -104 171 -88
rect -125 -181 -109 -147
rect 109 -181 125 -147
rect -285 -249 -251 -187
rect 251 -249 285 -187
rect -285 -283 -189 -249
rect 189 -283 285 -249
<< viali >>
rect -109 147 109 181
rect -171 -88 -137 88
rect 137 -88 171 88
rect -109 -181 109 -147
<< metal1 >>
rect -121 181 121 187
rect -121 147 -109 181
rect 109 147 121 181
rect -121 141 121 147
rect -177 88 -131 100
rect -177 -88 -171 88
rect -137 -88 -131 88
rect -177 -100 -131 -88
rect 131 88 177 100
rect 131 -88 137 88
rect 171 -88 177 88
rect 131 -100 177 -88
rect -121 -147 121 -141
rect -121 -181 -109 -147
rect 109 -181 121 -147
rect -121 -187 121 -181
<< properties >>
string FIXED_BBOX -268 -266 268 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 1.25 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
