magic
tech sky130A
magscale 1 2
timestamp 1668293870
<< pwell >>
rect -937 -310 937 310
<< nmos >>
rect -741 -100 -491 100
rect -433 -100 -183 100
rect -125 -100 125 100
rect 183 -100 433 100
rect 491 -100 741 100
<< ndiff >>
rect -799 88 -741 100
rect -799 -88 -787 88
rect -753 -88 -741 88
rect -799 -100 -741 -88
rect -491 88 -433 100
rect -491 -88 -479 88
rect -445 -88 -433 88
rect -491 -100 -433 -88
rect -183 88 -125 100
rect -183 -88 -171 88
rect -137 -88 -125 88
rect -183 -100 -125 -88
rect 125 88 183 100
rect 125 -88 137 88
rect 171 -88 183 88
rect 125 -100 183 -88
rect 433 88 491 100
rect 433 -88 445 88
rect 479 -88 491 88
rect 433 -100 491 -88
rect 741 88 799 100
rect 741 -88 753 88
rect 787 -88 799 88
rect 741 -100 799 -88
<< ndiffc >>
rect -787 -88 -753 88
rect -479 -88 -445 88
rect -171 -88 -137 88
rect 137 -88 171 88
rect 445 -88 479 88
rect 753 -88 787 88
<< psubdiff >>
rect -901 240 -805 274
rect 805 240 901 274
rect -901 178 -867 240
rect 867 178 901 240
rect -901 -240 -867 -178
rect 867 -240 901 -178
rect -901 -274 -805 -240
rect 805 -274 901 -240
<< psubdiffcont >>
rect -805 240 805 274
rect -901 -178 -867 178
rect 867 -178 901 178
rect -805 -274 805 -240
<< poly >>
rect -741 172 -491 188
rect -741 138 -725 172
rect -507 138 -491 172
rect -741 100 -491 138
rect -433 172 -183 188
rect -433 138 -417 172
rect -199 138 -183 172
rect -433 100 -183 138
rect -125 172 125 188
rect -125 138 -109 172
rect 109 138 125 172
rect -125 100 125 138
rect 183 172 433 188
rect 183 138 199 172
rect 417 138 433 172
rect 183 100 433 138
rect 491 172 741 188
rect 491 138 507 172
rect 725 138 741 172
rect 491 100 741 138
rect -741 -138 -491 -100
rect -741 -172 -725 -138
rect -507 -172 -491 -138
rect -741 -188 -491 -172
rect -433 -138 -183 -100
rect -433 -172 -417 -138
rect -199 -172 -183 -138
rect -433 -188 -183 -172
rect -125 -138 125 -100
rect -125 -172 -109 -138
rect 109 -172 125 -138
rect -125 -188 125 -172
rect 183 -138 433 -100
rect 183 -172 199 -138
rect 417 -172 433 -138
rect 183 -188 433 -172
rect 491 -138 741 -100
rect 491 -172 507 -138
rect 725 -172 741 -138
rect 491 -188 741 -172
<< polycont >>
rect -725 138 -507 172
rect -417 138 -199 172
rect -109 138 109 172
rect 199 138 417 172
rect 507 138 725 172
rect -725 -172 -507 -138
rect -417 -172 -199 -138
rect -109 -172 109 -138
rect 199 -172 417 -138
rect 507 -172 725 -138
<< locali >>
rect -901 240 -805 274
rect 805 240 901 274
rect -901 178 -867 240
rect 867 178 901 240
rect -741 138 -725 172
rect -507 138 -491 172
rect -433 138 -417 172
rect -199 138 -183 172
rect -125 138 -109 172
rect 109 138 125 172
rect 183 138 199 172
rect 417 138 433 172
rect 491 138 507 172
rect 725 138 741 172
rect -787 88 -753 104
rect -787 -104 -753 -88
rect -479 88 -445 104
rect -479 -104 -445 -88
rect -171 88 -137 104
rect -171 -104 -137 -88
rect 137 88 171 104
rect 137 -104 171 -88
rect 445 88 479 104
rect 445 -104 479 -88
rect 753 88 787 104
rect 753 -104 787 -88
rect -741 -172 -725 -138
rect -507 -172 -491 -138
rect -433 -172 -417 -138
rect -199 -172 -183 -138
rect -125 -172 -109 -138
rect 109 -172 125 -138
rect 183 -172 199 -138
rect 417 -172 433 -138
rect 491 -172 507 -138
rect 725 -172 741 -138
rect -901 -240 -867 -178
rect 867 -240 901 -178
rect -901 -274 -805 -240
rect 805 -274 901 -240
<< viali >>
rect -725 138 -507 172
rect -417 138 -199 172
rect -109 138 109 172
rect 199 138 417 172
rect 507 138 725 172
rect -787 -88 -753 88
rect -479 -88 -445 88
rect -171 -88 -137 88
rect 137 -88 171 88
rect 445 -88 479 88
rect 753 -88 787 88
rect -725 -172 -507 -138
rect -417 -172 -199 -138
rect -109 -172 109 -138
rect 199 -172 417 -138
rect 507 -172 725 -138
<< metal1 >>
rect -737 172 -495 178
rect -737 138 -725 172
rect -507 138 -495 172
rect -737 132 -495 138
rect -429 172 -187 178
rect -429 138 -417 172
rect -199 138 -187 172
rect -429 132 -187 138
rect -121 172 121 178
rect -121 138 -109 172
rect 109 138 121 172
rect -121 132 121 138
rect 187 172 429 178
rect 187 138 199 172
rect 417 138 429 172
rect 187 132 429 138
rect 495 172 737 178
rect 495 138 507 172
rect 725 138 737 172
rect 495 132 737 138
rect -793 88 -747 100
rect -793 -88 -787 88
rect -753 -88 -747 88
rect -793 -100 -747 -88
rect -485 88 -439 100
rect -485 -88 -479 88
rect -445 -88 -439 88
rect -485 -100 -439 -88
rect -177 88 -131 100
rect -177 -88 -171 88
rect -137 -88 -131 88
rect -177 -100 -131 -88
rect 131 88 177 100
rect 131 -88 137 88
rect 171 -88 177 88
rect 131 -100 177 -88
rect 439 88 485 100
rect 439 -88 445 88
rect 479 -88 485 88
rect 439 -100 485 -88
rect 747 88 793 100
rect 747 -88 753 88
rect 787 -88 793 88
rect 747 -100 793 -88
rect -737 -138 -495 -132
rect -737 -172 -725 -138
rect -507 -172 -495 -138
rect -737 -178 -495 -172
rect -429 -138 -187 -132
rect -429 -172 -417 -138
rect -199 -172 -187 -138
rect -429 -178 -187 -172
rect -121 -138 121 -132
rect -121 -172 -109 -138
rect 109 -172 121 -138
rect -121 -178 121 -172
rect 187 -138 429 -132
rect 187 -172 199 -138
rect 417 -172 429 -138
rect 187 -178 429 -172
rect 495 -138 737 -132
rect 495 -172 507 -138
rect 725 -172 737 -138
rect 495 -178 737 -172
<< properties >>
string FIXED_BBOX -884 -257 884 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 1.25 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
