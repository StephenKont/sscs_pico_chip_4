magic
tech sky130A
magscale 1 2
timestamp 1666549282
<< metal3 >>
rect -5507 7790 -180 8197
rect 10 8169 5507 8197
rect -5507 2799 -172 7790
rect 10 2827 5423 8169
rect 5487 2827 5507 8169
rect 10 2799 5507 2827
rect -5507 -2699 -172 2699
rect 10 2671 5507 2699
rect 10 -2671 5423 2671
rect 5487 -2671 5507 2671
rect 10 -2699 5507 -2671
rect -5507 -8197 -172 -2799
rect 10 -2827 5507 -2799
rect 10 -8169 5423 -2827
rect 5487 -8169 5507 -2827
rect 10 -8197 5507 -8169
<< via3 >>
rect 5423 2827 5487 8169
rect 5423 -2671 5487 2671
rect 5423 -8169 5487 -2827
<< mimcap >>
rect -5407 8057 -209 8097
rect -5407 2939 -5367 8057
rect -249 2939 -209 8057
rect -5407 2899 -209 2939
rect 110 8057 5308 8097
rect 110 2939 150 8057
rect 5268 2939 5308 8057
rect 110 2899 5308 2939
rect -5407 2559 -209 2599
rect -5407 -2559 -5367 2559
rect -249 -2559 -209 2559
rect -5407 -2599 -209 -2559
rect 110 2559 5308 2599
rect 110 -2559 150 2559
rect 5268 -2559 5308 2559
rect 110 -2599 5308 -2559
rect -5407 -2939 -209 -2899
rect -5407 -8057 -5367 -2939
rect -249 -8057 -209 -2939
rect -5407 -8097 -209 -8057
rect 110 -2939 5308 -2899
rect 110 -8057 150 -2939
rect 5268 -8057 5308 -2939
rect 110 -8097 5308 -8057
<< mimcapcontact >>
rect -5367 2939 -249 8057
rect 150 2939 5268 8057
rect -5367 -2559 -249 2559
rect 150 -2559 5268 2559
rect -5367 -8057 -249 -2939
rect 150 -8057 5268 -2939
<< metal4 >>
rect -2860 8058 -2756 8247
rect -141 8185 -37 8247
rect -5368 8057 -248 8058
rect -5368 2939 -5367 8057
rect -249 2939 -248 8057
rect -5368 2938 -248 2939
rect -2860 2560 -2756 2938
rect -141 2811 -14 8185
rect 2657 8058 2761 8247
rect 5376 8185 5480 8247
rect 5376 8169 5503 8185
rect 149 8057 5269 8058
rect 149 2939 150 8057
rect 5268 2939 5269 8057
rect 149 2938 5269 2939
rect -141 2687 -37 2811
rect -5368 2559 -248 2560
rect -5368 -2559 -5367 2559
rect -249 -2559 -248 2559
rect -5368 -2560 -248 -2559
rect -2860 -2938 -2756 -2560
rect -141 -2687 -14 2687
rect 2657 2560 2761 2938
rect 5376 2827 5423 8169
rect 5487 2827 5503 8169
rect 5376 2811 5503 2827
rect 5376 2687 5480 2811
rect 5376 2671 5503 2687
rect 149 2559 5269 2560
rect 149 -2559 150 2559
rect 5268 -2559 5269 2559
rect 149 -2560 5269 -2559
rect -141 -2811 -37 -2687
rect -5368 -2939 -248 -2938
rect -5368 -8057 -5367 -2939
rect -249 -8057 -248 -2939
rect -5368 -8058 -248 -8057
rect -2860 -8247 -2756 -8058
rect -141 -8185 -14 -2811
rect 2657 -2938 2761 -2560
rect 5376 -2671 5423 2671
rect 5487 -2671 5503 2671
rect 5376 -2687 5503 -2671
rect 5376 -2811 5480 -2687
rect 5376 -2827 5503 -2811
rect 149 -2939 5269 -2938
rect 149 -8057 150 -2939
rect 5268 -8057 5269 -2939
rect 149 -8058 5269 -8057
rect -141 -8247 -37 -8185
rect 2657 -8247 2761 -8058
rect 5376 -8169 5423 -2827
rect 5487 -8169 5503 -2827
rect 5376 -8185 5503 -8169
rect 5376 -8247 5480 -8185
<< properties >>
string FIXED_BBOX 10 2799 5408 8197
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25.992 l 25.992 val 1.371k carea 2.00 cperi 0.19 nx 2 ny 3 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
