magic
tech sky130A
magscale 1 2
timestamp 1666639277
<< pwell >>
rect -6519 -658 6519 658
<< mvnmos >>
rect -6291 -400 -6191 400
rect -6133 -400 -6033 400
rect -5975 -400 -5875 400
rect -5817 -400 -5717 400
rect -5659 -400 -5559 400
rect -5501 -400 -5401 400
rect -5343 -400 -5243 400
rect -5185 -400 -5085 400
rect -5027 -400 -4927 400
rect -4869 -400 -4769 400
rect -4711 -400 -4611 400
rect -4553 -400 -4453 400
rect -4395 -400 -4295 400
rect -4237 -400 -4137 400
rect -4079 -400 -3979 400
rect -3921 -400 -3821 400
rect -3763 -400 -3663 400
rect -3605 -400 -3505 400
rect -3447 -400 -3347 400
rect -3289 -400 -3189 400
rect -3131 -400 -3031 400
rect -2973 -400 -2873 400
rect -2815 -400 -2715 400
rect -2657 -400 -2557 400
rect -2499 -400 -2399 400
rect -2341 -400 -2241 400
rect -2183 -400 -2083 400
rect -2025 -400 -1925 400
rect -1867 -400 -1767 400
rect -1709 -400 -1609 400
rect -1551 -400 -1451 400
rect -1393 -400 -1293 400
rect -1235 -400 -1135 400
rect -1077 -400 -977 400
rect -919 -400 -819 400
rect -761 -400 -661 400
rect -603 -400 -503 400
rect -445 -400 -345 400
rect -287 -400 -187 400
rect -129 -400 -29 400
rect 29 -400 129 400
rect 187 -400 287 400
rect 345 -400 445 400
rect 503 -400 603 400
rect 661 -400 761 400
rect 819 -400 919 400
rect 977 -400 1077 400
rect 1135 -400 1235 400
rect 1293 -400 1393 400
rect 1451 -400 1551 400
rect 1609 -400 1709 400
rect 1767 -400 1867 400
rect 1925 -400 2025 400
rect 2083 -400 2183 400
rect 2241 -400 2341 400
rect 2399 -400 2499 400
rect 2557 -400 2657 400
rect 2715 -400 2815 400
rect 2873 -400 2973 400
rect 3031 -400 3131 400
rect 3189 -400 3289 400
rect 3347 -400 3447 400
rect 3505 -400 3605 400
rect 3663 -400 3763 400
rect 3821 -400 3921 400
rect 3979 -400 4079 400
rect 4137 -400 4237 400
rect 4295 -400 4395 400
rect 4453 -400 4553 400
rect 4611 -400 4711 400
rect 4769 -400 4869 400
rect 4927 -400 5027 400
rect 5085 -400 5185 400
rect 5243 -400 5343 400
rect 5401 -400 5501 400
rect 5559 -400 5659 400
rect 5717 -400 5817 400
rect 5875 -400 5975 400
rect 6033 -400 6133 400
rect 6191 -400 6291 400
<< mvndiff >>
rect -6349 388 -6291 400
rect -6349 -388 -6337 388
rect -6303 -388 -6291 388
rect -6349 -400 -6291 -388
rect -6191 388 -6133 400
rect -6191 -388 -6179 388
rect -6145 -388 -6133 388
rect -6191 -400 -6133 -388
rect -6033 388 -5975 400
rect -6033 -388 -6021 388
rect -5987 -388 -5975 388
rect -6033 -400 -5975 -388
rect -5875 388 -5817 400
rect -5875 -388 -5863 388
rect -5829 -388 -5817 388
rect -5875 -400 -5817 -388
rect -5717 388 -5659 400
rect -5717 -388 -5705 388
rect -5671 -388 -5659 388
rect -5717 -400 -5659 -388
rect -5559 388 -5501 400
rect -5559 -388 -5547 388
rect -5513 -388 -5501 388
rect -5559 -400 -5501 -388
rect -5401 388 -5343 400
rect -5401 -388 -5389 388
rect -5355 -388 -5343 388
rect -5401 -400 -5343 -388
rect -5243 388 -5185 400
rect -5243 -388 -5231 388
rect -5197 -388 -5185 388
rect -5243 -400 -5185 -388
rect -5085 388 -5027 400
rect -5085 -388 -5073 388
rect -5039 -388 -5027 388
rect -5085 -400 -5027 -388
rect -4927 388 -4869 400
rect -4927 -388 -4915 388
rect -4881 -388 -4869 388
rect -4927 -400 -4869 -388
rect -4769 388 -4711 400
rect -4769 -388 -4757 388
rect -4723 -388 -4711 388
rect -4769 -400 -4711 -388
rect -4611 388 -4553 400
rect -4611 -388 -4599 388
rect -4565 -388 -4553 388
rect -4611 -400 -4553 -388
rect -4453 388 -4395 400
rect -4453 -388 -4441 388
rect -4407 -388 -4395 388
rect -4453 -400 -4395 -388
rect -4295 388 -4237 400
rect -4295 -388 -4283 388
rect -4249 -388 -4237 388
rect -4295 -400 -4237 -388
rect -4137 388 -4079 400
rect -4137 -388 -4125 388
rect -4091 -388 -4079 388
rect -4137 -400 -4079 -388
rect -3979 388 -3921 400
rect -3979 -388 -3967 388
rect -3933 -388 -3921 388
rect -3979 -400 -3921 -388
rect -3821 388 -3763 400
rect -3821 -388 -3809 388
rect -3775 -388 -3763 388
rect -3821 -400 -3763 -388
rect -3663 388 -3605 400
rect -3663 -388 -3651 388
rect -3617 -388 -3605 388
rect -3663 -400 -3605 -388
rect -3505 388 -3447 400
rect -3505 -388 -3493 388
rect -3459 -388 -3447 388
rect -3505 -400 -3447 -388
rect -3347 388 -3289 400
rect -3347 -388 -3335 388
rect -3301 -388 -3289 388
rect -3347 -400 -3289 -388
rect -3189 388 -3131 400
rect -3189 -388 -3177 388
rect -3143 -388 -3131 388
rect -3189 -400 -3131 -388
rect -3031 388 -2973 400
rect -3031 -388 -3019 388
rect -2985 -388 -2973 388
rect -3031 -400 -2973 -388
rect -2873 388 -2815 400
rect -2873 -388 -2861 388
rect -2827 -388 -2815 388
rect -2873 -400 -2815 -388
rect -2715 388 -2657 400
rect -2715 -388 -2703 388
rect -2669 -388 -2657 388
rect -2715 -400 -2657 -388
rect -2557 388 -2499 400
rect -2557 -388 -2545 388
rect -2511 -388 -2499 388
rect -2557 -400 -2499 -388
rect -2399 388 -2341 400
rect -2399 -388 -2387 388
rect -2353 -388 -2341 388
rect -2399 -400 -2341 -388
rect -2241 388 -2183 400
rect -2241 -388 -2229 388
rect -2195 -388 -2183 388
rect -2241 -400 -2183 -388
rect -2083 388 -2025 400
rect -2083 -388 -2071 388
rect -2037 -388 -2025 388
rect -2083 -400 -2025 -388
rect -1925 388 -1867 400
rect -1925 -388 -1913 388
rect -1879 -388 -1867 388
rect -1925 -400 -1867 -388
rect -1767 388 -1709 400
rect -1767 -388 -1755 388
rect -1721 -388 -1709 388
rect -1767 -400 -1709 -388
rect -1609 388 -1551 400
rect -1609 -388 -1597 388
rect -1563 -388 -1551 388
rect -1609 -400 -1551 -388
rect -1451 388 -1393 400
rect -1451 -388 -1439 388
rect -1405 -388 -1393 388
rect -1451 -400 -1393 -388
rect -1293 388 -1235 400
rect -1293 -388 -1281 388
rect -1247 -388 -1235 388
rect -1293 -400 -1235 -388
rect -1135 388 -1077 400
rect -1135 -388 -1123 388
rect -1089 -388 -1077 388
rect -1135 -400 -1077 -388
rect -977 388 -919 400
rect -977 -388 -965 388
rect -931 -388 -919 388
rect -977 -400 -919 -388
rect -819 388 -761 400
rect -819 -388 -807 388
rect -773 -388 -761 388
rect -819 -400 -761 -388
rect -661 388 -603 400
rect -661 -388 -649 388
rect -615 -388 -603 388
rect -661 -400 -603 -388
rect -503 388 -445 400
rect -503 -388 -491 388
rect -457 -388 -445 388
rect -503 -400 -445 -388
rect -345 388 -287 400
rect -345 -388 -333 388
rect -299 -388 -287 388
rect -345 -400 -287 -388
rect -187 388 -129 400
rect -187 -388 -175 388
rect -141 -388 -129 388
rect -187 -400 -129 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 129 388 187 400
rect 129 -388 141 388
rect 175 -388 187 388
rect 129 -400 187 -388
rect 287 388 345 400
rect 287 -388 299 388
rect 333 -388 345 388
rect 287 -400 345 -388
rect 445 388 503 400
rect 445 -388 457 388
rect 491 -388 503 388
rect 445 -400 503 -388
rect 603 388 661 400
rect 603 -388 615 388
rect 649 -388 661 388
rect 603 -400 661 -388
rect 761 388 819 400
rect 761 -388 773 388
rect 807 -388 819 388
rect 761 -400 819 -388
rect 919 388 977 400
rect 919 -388 931 388
rect 965 -388 977 388
rect 919 -400 977 -388
rect 1077 388 1135 400
rect 1077 -388 1089 388
rect 1123 -388 1135 388
rect 1077 -400 1135 -388
rect 1235 388 1293 400
rect 1235 -388 1247 388
rect 1281 -388 1293 388
rect 1235 -400 1293 -388
rect 1393 388 1451 400
rect 1393 -388 1405 388
rect 1439 -388 1451 388
rect 1393 -400 1451 -388
rect 1551 388 1609 400
rect 1551 -388 1563 388
rect 1597 -388 1609 388
rect 1551 -400 1609 -388
rect 1709 388 1767 400
rect 1709 -388 1721 388
rect 1755 -388 1767 388
rect 1709 -400 1767 -388
rect 1867 388 1925 400
rect 1867 -388 1879 388
rect 1913 -388 1925 388
rect 1867 -400 1925 -388
rect 2025 388 2083 400
rect 2025 -388 2037 388
rect 2071 -388 2083 388
rect 2025 -400 2083 -388
rect 2183 388 2241 400
rect 2183 -388 2195 388
rect 2229 -388 2241 388
rect 2183 -400 2241 -388
rect 2341 388 2399 400
rect 2341 -388 2353 388
rect 2387 -388 2399 388
rect 2341 -400 2399 -388
rect 2499 388 2557 400
rect 2499 -388 2511 388
rect 2545 -388 2557 388
rect 2499 -400 2557 -388
rect 2657 388 2715 400
rect 2657 -388 2669 388
rect 2703 -388 2715 388
rect 2657 -400 2715 -388
rect 2815 388 2873 400
rect 2815 -388 2827 388
rect 2861 -388 2873 388
rect 2815 -400 2873 -388
rect 2973 388 3031 400
rect 2973 -388 2985 388
rect 3019 -388 3031 388
rect 2973 -400 3031 -388
rect 3131 388 3189 400
rect 3131 -388 3143 388
rect 3177 -388 3189 388
rect 3131 -400 3189 -388
rect 3289 388 3347 400
rect 3289 -388 3301 388
rect 3335 -388 3347 388
rect 3289 -400 3347 -388
rect 3447 388 3505 400
rect 3447 -388 3459 388
rect 3493 -388 3505 388
rect 3447 -400 3505 -388
rect 3605 388 3663 400
rect 3605 -388 3617 388
rect 3651 -388 3663 388
rect 3605 -400 3663 -388
rect 3763 388 3821 400
rect 3763 -388 3775 388
rect 3809 -388 3821 388
rect 3763 -400 3821 -388
rect 3921 388 3979 400
rect 3921 -388 3933 388
rect 3967 -388 3979 388
rect 3921 -400 3979 -388
rect 4079 388 4137 400
rect 4079 -388 4091 388
rect 4125 -388 4137 388
rect 4079 -400 4137 -388
rect 4237 388 4295 400
rect 4237 -388 4249 388
rect 4283 -388 4295 388
rect 4237 -400 4295 -388
rect 4395 388 4453 400
rect 4395 -388 4407 388
rect 4441 -388 4453 388
rect 4395 -400 4453 -388
rect 4553 388 4611 400
rect 4553 -388 4565 388
rect 4599 -388 4611 388
rect 4553 -400 4611 -388
rect 4711 388 4769 400
rect 4711 -388 4723 388
rect 4757 -388 4769 388
rect 4711 -400 4769 -388
rect 4869 388 4927 400
rect 4869 -388 4881 388
rect 4915 -388 4927 388
rect 4869 -400 4927 -388
rect 5027 388 5085 400
rect 5027 -388 5039 388
rect 5073 -388 5085 388
rect 5027 -400 5085 -388
rect 5185 388 5243 400
rect 5185 -388 5197 388
rect 5231 -388 5243 388
rect 5185 -400 5243 -388
rect 5343 388 5401 400
rect 5343 -388 5355 388
rect 5389 -388 5401 388
rect 5343 -400 5401 -388
rect 5501 388 5559 400
rect 5501 -388 5513 388
rect 5547 -388 5559 388
rect 5501 -400 5559 -388
rect 5659 388 5717 400
rect 5659 -388 5671 388
rect 5705 -388 5717 388
rect 5659 -400 5717 -388
rect 5817 388 5875 400
rect 5817 -388 5829 388
rect 5863 -388 5875 388
rect 5817 -400 5875 -388
rect 5975 388 6033 400
rect 5975 -388 5987 388
rect 6021 -388 6033 388
rect 5975 -400 6033 -388
rect 6133 388 6191 400
rect 6133 -388 6145 388
rect 6179 -388 6191 388
rect 6133 -400 6191 -388
rect 6291 388 6349 400
rect 6291 -388 6303 388
rect 6337 -388 6349 388
rect 6291 -400 6349 -388
<< mvndiffc >>
rect -6337 -388 -6303 388
rect -6179 -388 -6145 388
rect -6021 -388 -5987 388
rect -5863 -388 -5829 388
rect -5705 -388 -5671 388
rect -5547 -388 -5513 388
rect -5389 -388 -5355 388
rect -5231 -388 -5197 388
rect -5073 -388 -5039 388
rect -4915 -388 -4881 388
rect -4757 -388 -4723 388
rect -4599 -388 -4565 388
rect -4441 -388 -4407 388
rect -4283 -388 -4249 388
rect -4125 -388 -4091 388
rect -3967 -388 -3933 388
rect -3809 -388 -3775 388
rect -3651 -388 -3617 388
rect -3493 -388 -3459 388
rect -3335 -388 -3301 388
rect -3177 -388 -3143 388
rect -3019 -388 -2985 388
rect -2861 -388 -2827 388
rect -2703 -388 -2669 388
rect -2545 -388 -2511 388
rect -2387 -388 -2353 388
rect -2229 -388 -2195 388
rect -2071 -388 -2037 388
rect -1913 -388 -1879 388
rect -1755 -388 -1721 388
rect -1597 -388 -1563 388
rect -1439 -388 -1405 388
rect -1281 -388 -1247 388
rect -1123 -388 -1089 388
rect -965 -388 -931 388
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
rect 931 -388 965 388
rect 1089 -388 1123 388
rect 1247 -388 1281 388
rect 1405 -388 1439 388
rect 1563 -388 1597 388
rect 1721 -388 1755 388
rect 1879 -388 1913 388
rect 2037 -388 2071 388
rect 2195 -388 2229 388
rect 2353 -388 2387 388
rect 2511 -388 2545 388
rect 2669 -388 2703 388
rect 2827 -388 2861 388
rect 2985 -388 3019 388
rect 3143 -388 3177 388
rect 3301 -388 3335 388
rect 3459 -388 3493 388
rect 3617 -388 3651 388
rect 3775 -388 3809 388
rect 3933 -388 3967 388
rect 4091 -388 4125 388
rect 4249 -388 4283 388
rect 4407 -388 4441 388
rect 4565 -388 4599 388
rect 4723 -388 4757 388
rect 4881 -388 4915 388
rect 5039 -388 5073 388
rect 5197 -388 5231 388
rect 5355 -388 5389 388
rect 5513 -388 5547 388
rect 5671 -388 5705 388
rect 5829 -388 5863 388
rect 5987 -388 6021 388
rect 6145 -388 6179 388
rect 6303 -388 6337 388
<< mvpsubdiff >>
rect -6483 610 6483 622
rect -6483 576 -6375 610
rect 6375 576 6483 610
rect -6483 564 6483 576
rect -6483 514 -6425 564
rect -6483 -514 -6471 514
rect -6437 -514 -6425 514
rect 6425 514 6483 564
rect -6483 -564 -6425 -514
rect 6425 -514 6437 514
rect 6471 -514 6483 514
rect 6425 -564 6483 -514
rect -6483 -576 6483 -564
rect -6483 -610 -6375 -576
rect 6375 -610 6483 -576
rect -6483 -622 6483 -610
<< mvpsubdiffcont >>
rect -6375 576 6375 610
rect -6471 -514 -6437 514
rect 6437 -514 6471 514
rect -6375 -610 6375 -576
<< poly >>
rect -6291 472 -6191 488
rect -6291 438 -6275 472
rect -6207 438 -6191 472
rect -6291 400 -6191 438
rect -6133 472 -6033 488
rect -6133 438 -6117 472
rect -6049 438 -6033 472
rect -6133 400 -6033 438
rect -5975 472 -5875 488
rect -5975 438 -5959 472
rect -5891 438 -5875 472
rect -5975 400 -5875 438
rect -5817 472 -5717 488
rect -5817 438 -5801 472
rect -5733 438 -5717 472
rect -5817 400 -5717 438
rect -5659 472 -5559 488
rect -5659 438 -5643 472
rect -5575 438 -5559 472
rect -5659 400 -5559 438
rect -5501 472 -5401 488
rect -5501 438 -5485 472
rect -5417 438 -5401 472
rect -5501 400 -5401 438
rect -5343 472 -5243 488
rect -5343 438 -5327 472
rect -5259 438 -5243 472
rect -5343 400 -5243 438
rect -5185 472 -5085 488
rect -5185 438 -5169 472
rect -5101 438 -5085 472
rect -5185 400 -5085 438
rect -5027 472 -4927 488
rect -5027 438 -5011 472
rect -4943 438 -4927 472
rect -5027 400 -4927 438
rect -4869 472 -4769 488
rect -4869 438 -4853 472
rect -4785 438 -4769 472
rect -4869 400 -4769 438
rect -4711 472 -4611 488
rect -4711 438 -4695 472
rect -4627 438 -4611 472
rect -4711 400 -4611 438
rect -4553 472 -4453 488
rect -4553 438 -4537 472
rect -4469 438 -4453 472
rect -4553 400 -4453 438
rect -4395 472 -4295 488
rect -4395 438 -4379 472
rect -4311 438 -4295 472
rect -4395 400 -4295 438
rect -4237 472 -4137 488
rect -4237 438 -4221 472
rect -4153 438 -4137 472
rect -4237 400 -4137 438
rect -4079 472 -3979 488
rect -4079 438 -4063 472
rect -3995 438 -3979 472
rect -4079 400 -3979 438
rect -3921 472 -3821 488
rect -3921 438 -3905 472
rect -3837 438 -3821 472
rect -3921 400 -3821 438
rect -3763 472 -3663 488
rect -3763 438 -3747 472
rect -3679 438 -3663 472
rect -3763 400 -3663 438
rect -3605 472 -3505 488
rect -3605 438 -3589 472
rect -3521 438 -3505 472
rect -3605 400 -3505 438
rect -3447 472 -3347 488
rect -3447 438 -3431 472
rect -3363 438 -3347 472
rect -3447 400 -3347 438
rect -3289 472 -3189 488
rect -3289 438 -3273 472
rect -3205 438 -3189 472
rect -3289 400 -3189 438
rect -3131 472 -3031 488
rect -3131 438 -3115 472
rect -3047 438 -3031 472
rect -3131 400 -3031 438
rect -2973 472 -2873 488
rect -2973 438 -2957 472
rect -2889 438 -2873 472
rect -2973 400 -2873 438
rect -2815 472 -2715 488
rect -2815 438 -2799 472
rect -2731 438 -2715 472
rect -2815 400 -2715 438
rect -2657 472 -2557 488
rect -2657 438 -2641 472
rect -2573 438 -2557 472
rect -2657 400 -2557 438
rect -2499 472 -2399 488
rect -2499 438 -2483 472
rect -2415 438 -2399 472
rect -2499 400 -2399 438
rect -2341 472 -2241 488
rect -2341 438 -2325 472
rect -2257 438 -2241 472
rect -2341 400 -2241 438
rect -2183 472 -2083 488
rect -2183 438 -2167 472
rect -2099 438 -2083 472
rect -2183 400 -2083 438
rect -2025 472 -1925 488
rect -2025 438 -2009 472
rect -1941 438 -1925 472
rect -2025 400 -1925 438
rect -1867 472 -1767 488
rect -1867 438 -1851 472
rect -1783 438 -1767 472
rect -1867 400 -1767 438
rect -1709 472 -1609 488
rect -1709 438 -1693 472
rect -1625 438 -1609 472
rect -1709 400 -1609 438
rect -1551 472 -1451 488
rect -1551 438 -1535 472
rect -1467 438 -1451 472
rect -1551 400 -1451 438
rect -1393 472 -1293 488
rect -1393 438 -1377 472
rect -1309 438 -1293 472
rect -1393 400 -1293 438
rect -1235 472 -1135 488
rect -1235 438 -1219 472
rect -1151 438 -1135 472
rect -1235 400 -1135 438
rect -1077 472 -977 488
rect -1077 438 -1061 472
rect -993 438 -977 472
rect -1077 400 -977 438
rect -919 472 -819 488
rect -919 438 -903 472
rect -835 438 -819 472
rect -919 400 -819 438
rect -761 472 -661 488
rect -761 438 -745 472
rect -677 438 -661 472
rect -761 400 -661 438
rect -603 472 -503 488
rect -603 438 -587 472
rect -519 438 -503 472
rect -603 400 -503 438
rect -445 472 -345 488
rect -445 438 -429 472
rect -361 438 -345 472
rect -445 400 -345 438
rect -287 472 -187 488
rect -287 438 -271 472
rect -203 438 -187 472
rect -287 400 -187 438
rect -129 472 -29 488
rect -129 438 -113 472
rect -45 438 -29 472
rect -129 400 -29 438
rect 29 472 129 488
rect 29 438 45 472
rect 113 438 129 472
rect 29 400 129 438
rect 187 472 287 488
rect 187 438 203 472
rect 271 438 287 472
rect 187 400 287 438
rect 345 472 445 488
rect 345 438 361 472
rect 429 438 445 472
rect 345 400 445 438
rect 503 472 603 488
rect 503 438 519 472
rect 587 438 603 472
rect 503 400 603 438
rect 661 472 761 488
rect 661 438 677 472
rect 745 438 761 472
rect 661 400 761 438
rect 819 472 919 488
rect 819 438 835 472
rect 903 438 919 472
rect 819 400 919 438
rect 977 472 1077 488
rect 977 438 993 472
rect 1061 438 1077 472
rect 977 400 1077 438
rect 1135 472 1235 488
rect 1135 438 1151 472
rect 1219 438 1235 472
rect 1135 400 1235 438
rect 1293 472 1393 488
rect 1293 438 1309 472
rect 1377 438 1393 472
rect 1293 400 1393 438
rect 1451 472 1551 488
rect 1451 438 1467 472
rect 1535 438 1551 472
rect 1451 400 1551 438
rect 1609 472 1709 488
rect 1609 438 1625 472
rect 1693 438 1709 472
rect 1609 400 1709 438
rect 1767 472 1867 488
rect 1767 438 1783 472
rect 1851 438 1867 472
rect 1767 400 1867 438
rect 1925 472 2025 488
rect 1925 438 1941 472
rect 2009 438 2025 472
rect 1925 400 2025 438
rect 2083 472 2183 488
rect 2083 438 2099 472
rect 2167 438 2183 472
rect 2083 400 2183 438
rect 2241 472 2341 488
rect 2241 438 2257 472
rect 2325 438 2341 472
rect 2241 400 2341 438
rect 2399 472 2499 488
rect 2399 438 2415 472
rect 2483 438 2499 472
rect 2399 400 2499 438
rect 2557 472 2657 488
rect 2557 438 2573 472
rect 2641 438 2657 472
rect 2557 400 2657 438
rect 2715 472 2815 488
rect 2715 438 2731 472
rect 2799 438 2815 472
rect 2715 400 2815 438
rect 2873 472 2973 488
rect 2873 438 2889 472
rect 2957 438 2973 472
rect 2873 400 2973 438
rect 3031 472 3131 488
rect 3031 438 3047 472
rect 3115 438 3131 472
rect 3031 400 3131 438
rect 3189 472 3289 488
rect 3189 438 3205 472
rect 3273 438 3289 472
rect 3189 400 3289 438
rect 3347 472 3447 488
rect 3347 438 3363 472
rect 3431 438 3447 472
rect 3347 400 3447 438
rect 3505 472 3605 488
rect 3505 438 3521 472
rect 3589 438 3605 472
rect 3505 400 3605 438
rect 3663 472 3763 488
rect 3663 438 3679 472
rect 3747 438 3763 472
rect 3663 400 3763 438
rect 3821 472 3921 488
rect 3821 438 3837 472
rect 3905 438 3921 472
rect 3821 400 3921 438
rect 3979 472 4079 488
rect 3979 438 3995 472
rect 4063 438 4079 472
rect 3979 400 4079 438
rect 4137 472 4237 488
rect 4137 438 4153 472
rect 4221 438 4237 472
rect 4137 400 4237 438
rect 4295 472 4395 488
rect 4295 438 4311 472
rect 4379 438 4395 472
rect 4295 400 4395 438
rect 4453 472 4553 488
rect 4453 438 4469 472
rect 4537 438 4553 472
rect 4453 400 4553 438
rect 4611 472 4711 488
rect 4611 438 4627 472
rect 4695 438 4711 472
rect 4611 400 4711 438
rect 4769 472 4869 488
rect 4769 438 4785 472
rect 4853 438 4869 472
rect 4769 400 4869 438
rect 4927 472 5027 488
rect 4927 438 4943 472
rect 5011 438 5027 472
rect 4927 400 5027 438
rect 5085 472 5185 488
rect 5085 438 5101 472
rect 5169 438 5185 472
rect 5085 400 5185 438
rect 5243 472 5343 488
rect 5243 438 5259 472
rect 5327 438 5343 472
rect 5243 400 5343 438
rect 5401 472 5501 488
rect 5401 438 5417 472
rect 5485 438 5501 472
rect 5401 400 5501 438
rect 5559 472 5659 488
rect 5559 438 5575 472
rect 5643 438 5659 472
rect 5559 400 5659 438
rect 5717 472 5817 488
rect 5717 438 5733 472
rect 5801 438 5817 472
rect 5717 400 5817 438
rect 5875 472 5975 488
rect 5875 438 5891 472
rect 5959 438 5975 472
rect 5875 400 5975 438
rect 6033 472 6133 488
rect 6033 438 6049 472
rect 6117 438 6133 472
rect 6033 400 6133 438
rect 6191 472 6291 488
rect 6191 438 6207 472
rect 6275 438 6291 472
rect 6191 400 6291 438
rect -6291 -438 -6191 -400
rect -6291 -472 -6275 -438
rect -6207 -472 -6191 -438
rect -6291 -488 -6191 -472
rect -6133 -438 -6033 -400
rect -6133 -472 -6117 -438
rect -6049 -472 -6033 -438
rect -6133 -488 -6033 -472
rect -5975 -438 -5875 -400
rect -5975 -472 -5959 -438
rect -5891 -472 -5875 -438
rect -5975 -488 -5875 -472
rect -5817 -438 -5717 -400
rect -5817 -472 -5801 -438
rect -5733 -472 -5717 -438
rect -5817 -488 -5717 -472
rect -5659 -438 -5559 -400
rect -5659 -472 -5643 -438
rect -5575 -472 -5559 -438
rect -5659 -488 -5559 -472
rect -5501 -438 -5401 -400
rect -5501 -472 -5485 -438
rect -5417 -472 -5401 -438
rect -5501 -488 -5401 -472
rect -5343 -438 -5243 -400
rect -5343 -472 -5327 -438
rect -5259 -472 -5243 -438
rect -5343 -488 -5243 -472
rect -5185 -438 -5085 -400
rect -5185 -472 -5169 -438
rect -5101 -472 -5085 -438
rect -5185 -488 -5085 -472
rect -5027 -438 -4927 -400
rect -5027 -472 -5011 -438
rect -4943 -472 -4927 -438
rect -5027 -488 -4927 -472
rect -4869 -438 -4769 -400
rect -4869 -472 -4853 -438
rect -4785 -472 -4769 -438
rect -4869 -488 -4769 -472
rect -4711 -438 -4611 -400
rect -4711 -472 -4695 -438
rect -4627 -472 -4611 -438
rect -4711 -488 -4611 -472
rect -4553 -438 -4453 -400
rect -4553 -472 -4537 -438
rect -4469 -472 -4453 -438
rect -4553 -488 -4453 -472
rect -4395 -438 -4295 -400
rect -4395 -472 -4379 -438
rect -4311 -472 -4295 -438
rect -4395 -488 -4295 -472
rect -4237 -438 -4137 -400
rect -4237 -472 -4221 -438
rect -4153 -472 -4137 -438
rect -4237 -488 -4137 -472
rect -4079 -438 -3979 -400
rect -4079 -472 -4063 -438
rect -3995 -472 -3979 -438
rect -4079 -488 -3979 -472
rect -3921 -438 -3821 -400
rect -3921 -472 -3905 -438
rect -3837 -472 -3821 -438
rect -3921 -488 -3821 -472
rect -3763 -438 -3663 -400
rect -3763 -472 -3747 -438
rect -3679 -472 -3663 -438
rect -3763 -488 -3663 -472
rect -3605 -438 -3505 -400
rect -3605 -472 -3589 -438
rect -3521 -472 -3505 -438
rect -3605 -488 -3505 -472
rect -3447 -438 -3347 -400
rect -3447 -472 -3431 -438
rect -3363 -472 -3347 -438
rect -3447 -488 -3347 -472
rect -3289 -438 -3189 -400
rect -3289 -472 -3273 -438
rect -3205 -472 -3189 -438
rect -3289 -488 -3189 -472
rect -3131 -438 -3031 -400
rect -3131 -472 -3115 -438
rect -3047 -472 -3031 -438
rect -3131 -488 -3031 -472
rect -2973 -438 -2873 -400
rect -2973 -472 -2957 -438
rect -2889 -472 -2873 -438
rect -2973 -488 -2873 -472
rect -2815 -438 -2715 -400
rect -2815 -472 -2799 -438
rect -2731 -472 -2715 -438
rect -2815 -488 -2715 -472
rect -2657 -438 -2557 -400
rect -2657 -472 -2641 -438
rect -2573 -472 -2557 -438
rect -2657 -488 -2557 -472
rect -2499 -438 -2399 -400
rect -2499 -472 -2483 -438
rect -2415 -472 -2399 -438
rect -2499 -488 -2399 -472
rect -2341 -438 -2241 -400
rect -2341 -472 -2325 -438
rect -2257 -472 -2241 -438
rect -2341 -488 -2241 -472
rect -2183 -438 -2083 -400
rect -2183 -472 -2167 -438
rect -2099 -472 -2083 -438
rect -2183 -488 -2083 -472
rect -2025 -438 -1925 -400
rect -2025 -472 -2009 -438
rect -1941 -472 -1925 -438
rect -2025 -488 -1925 -472
rect -1867 -438 -1767 -400
rect -1867 -472 -1851 -438
rect -1783 -472 -1767 -438
rect -1867 -488 -1767 -472
rect -1709 -438 -1609 -400
rect -1709 -472 -1693 -438
rect -1625 -472 -1609 -438
rect -1709 -488 -1609 -472
rect -1551 -438 -1451 -400
rect -1551 -472 -1535 -438
rect -1467 -472 -1451 -438
rect -1551 -488 -1451 -472
rect -1393 -438 -1293 -400
rect -1393 -472 -1377 -438
rect -1309 -472 -1293 -438
rect -1393 -488 -1293 -472
rect -1235 -438 -1135 -400
rect -1235 -472 -1219 -438
rect -1151 -472 -1135 -438
rect -1235 -488 -1135 -472
rect -1077 -438 -977 -400
rect -1077 -472 -1061 -438
rect -993 -472 -977 -438
rect -1077 -488 -977 -472
rect -919 -438 -819 -400
rect -919 -472 -903 -438
rect -835 -472 -819 -438
rect -919 -488 -819 -472
rect -761 -438 -661 -400
rect -761 -472 -745 -438
rect -677 -472 -661 -438
rect -761 -488 -661 -472
rect -603 -438 -503 -400
rect -603 -472 -587 -438
rect -519 -472 -503 -438
rect -603 -488 -503 -472
rect -445 -438 -345 -400
rect -445 -472 -429 -438
rect -361 -472 -345 -438
rect -445 -488 -345 -472
rect -287 -438 -187 -400
rect -287 -472 -271 -438
rect -203 -472 -187 -438
rect -287 -488 -187 -472
rect -129 -438 -29 -400
rect -129 -472 -113 -438
rect -45 -472 -29 -438
rect -129 -488 -29 -472
rect 29 -438 129 -400
rect 29 -472 45 -438
rect 113 -472 129 -438
rect 29 -488 129 -472
rect 187 -438 287 -400
rect 187 -472 203 -438
rect 271 -472 287 -438
rect 187 -488 287 -472
rect 345 -438 445 -400
rect 345 -472 361 -438
rect 429 -472 445 -438
rect 345 -488 445 -472
rect 503 -438 603 -400
rect 503 -472 519 -438
rect 587 -472 603 -438
rect 503 -488 603 -472
rect 661 -438 761 -400
rect 661 -472 677 -438
rect 745 -472 761 -438
rect 661 -488 761 -472
rect 819 -438 919 -400
rect 819 -472 835 -438
rect 903 -472 919 -438
rect 819 -488 919 -472
rect 977 -438 1077 -400
rect 977 -472 993 -438
rect 1061 -472 1077 -438
rect 977 -488 1077 -472
rect 1135 -438 1235 -400
rect 1135 -472 1151 -438
rect 1219 -472 1235 -438
rect 1135 -488 1235 -472
rect 1293 -438 1393 -400
rect 1293 -472 1309 -438
rect 1377 -472 1393 -438
rect 1293 -488 1393 -472
rect 1451 -438 1551 -400
rect 1451 -472 1467 -438
rect 1535 -472 1551 -438
rect 1451 -488 1551 -472
rect 1609 -438 1709 -400
rect 1609 -472 1625 -438
rect 1693 -472 1709 -438
rect 1609 -488 1709 -472
rect 1767 -438 1867 -400
rect 1767 -472 1783 -438
rect 1851 -472 1867 -438
rect 1767 -488 1867 -472
rect 1925 -438 2025 -400
rect 1925 -472 1941 -438
rect 2009 -472 2025 -438
rect 1925 -488 2025 -472
rect 2083 -438 2183 -400
rect 2083 -472 2099 -438
rect 2167 -472 2183 -438
rect 2083 -488 2183 -472
rect 2241 -438 2341 -400
rect 2241 -472 2257 -438
rect 2325 -472 2341 -438
rect 2241 -488 2341 -472
rect 2399 -438 2499 -400
rect 2399 -472 2415 -438
rect 2483 -472 2499 -438
rect 2399 -488 2499 -472
rect 2557 -438 2657 -400
rect 2557 -472 2573 -438
rect 2641 -472 2657 -438
rect 2557 -488 2657 -472
rect 2715 -438 2815 -400
rect 2715 -472 2731 -438
rect 2799 -472 2815 -438
rect 2715 -488 2815 -472
rect 2873 -438 2973 -400
rect 2873 -472 2889 -438
rect 2957 -472 2973 -438
rect 2873 -488 2973 -472
rect 3031 -438 3131 -400
rect 3031 -472 3047 -438
rect 3115 -472 3131 -438
rect 3031 -488 3131 -472
rect 3189 -438 3289 -400
rect 3189 -472 3205 -438
rect 3273 -472 3289 -438
rect 3189 -488 3289 -472
rect 3347 -438 3447 -400
rect 3347 -472 3363 -438
rect 3431 -472 3447 -438
rect 3347 -488 3447 -472
rect 3505 -438 3605 -400
rect 3505 -472 3521 -438
rect 3589 -472 3605 -438
rect 3505 -488 3605 -472
rect 3663 -438 3763 -400
rect 3663 -472 3679 -438
rect 3747 -472 3763 -438
rect 3663 -488 3763 -472
rect 3821 -438 3921 -400
rect 3821 -472 3837 -438
rect 3905 -472 3921 -438
rect 3821 -488 3921 -472
rect 3979 -438 4079 -400
rect 3979 -472 3995 -438
rect 4063 -472 4079 -438
rect 3979 -488 4079 -472
rect 4137 -438 4237 -400
rect 4137 -472 4153 -438
rect 4221 -472 4237 -438
rect 4137 -488 4237 -472
rect 4295 -438 4395 -400
rect 4295 -472 4311 -438
rect 4379 -472 4395 -438
rect 4295 -488 4395 -472
rect 4453 -438 4553 -400
rect 4453 -472 4469 -438
rect 4537 -472 4553 -438
rect 4453 -488 4553 -472
rect 4611 -438 4711 -400
rect 4611 -472 4627 -438
rect 4695 -472 4711 -438
rect 4611 -488 4711 -472
rect 4769 -438 4869 -400
rect 4769 -472 4785 -438
rect 4853 -472 4869 -438
rect 4769 -488 4869 -472
rect 4927 -438 5027 -400
rect 4927 -472 4943 -438
rect 5011 -472 5027 -438
rect 4927 -488 5027 -472
rect 5085 -438 5185 -400
rect 5085 -472 5101 -438
rect 5169 -472 5185 -438
rect 5085 -488 5185 -472
rect 5243 -438 5343 -400
rect 5243 -472 5259 -438
rect 5327 -472 5343 -438
rect 5243 -488 5343 -472
rect 5401 -438 5501 -400
rect 5401 -472 5417 -438
rect 5485 -472 5501 -438
rect 5401 -488 5501 -472
rect 5559 -438 5659 -400
rect 5559 -472 5575 -438
rect 5643 -472 5659 -438
rect 5559 -488 5659 -472
rect 5717 -438 5817 -400
rect 5717 -472 5733 -438
rect 5801 -472 5817 -438
rect 5717 -488 5817 -472
rect 5875 -438 5975 -400
rect 5875 -472 5891 -438
rect 5959 -472 5975 -438
rect 5875 -488 5975 -472
rect 6033 -438 6133 -400
rect 6033 -472 6049 -438
rect 6117 -472 6133 -438
rect 6033 -488 6133 -472
rect 6191 -438 6291 -400
rect 6191 -472 6207 -438
rect 6275 -472 6291 -438
rect 6191 -488 6291 -472
<< polycont >>
rect -6275 438 -6207 472
rect -6117 438 -6049 472
rect -5959 438 -5891 472
rect -5801 438 -5733 472
rect -5643 438 -5575 472
rect -5485 438 -5417 472
rect -5327 438 -5259 472
rect -5169 438 -5101 472
rect -5011 438 -4943 472
rect -4853 438 -4785 472
rect -4695 438 -4627 472
rect -4537 438 -4469 472
rect -4379 438 -4311 472
rect -4221 438 -4153 472
rect -4063 438 -3995 472
rect -3905 438 -3837 472
rect -3747 438 -3679 472
rect -3589 438 -3521 472
rect -3431 438 -3363 472
rect -3273 438 -3205 472
rect -3115 438 -3047 472
rect -2957 438 -2889 472
rect -2799 438 -2731 472
rect -2641 438 -2573 472
rect -2483 438 -2415 472
rect -2325 438 -2257 472
rect -2167 438 -2099 472
rect -2009 438 -1941 472
rect -1851 438 -1783 472
rect -1693 438 -1625 472
rect -1535 438 -1467 472
rect -1377 438 -1309 472
rect -1219 438 -1151 472
rect -1061 438 -993 472
rect -903 438 -835 472
rect -745 438 -677 472
rect -587 438 -519 472
rect -429 438 -361 472
rect -271 438 -203 472
rect -113 438 -45 472
rect 45 438 113 472
rect 203 438 271 472
rect 361 438 429 472
rect 519 438 587 472
rect 677 438 745 472
rect 835 438 903 472
rect 993 438 1061 472
rect 1151 438 1219 472
rect 1309 438 1377 472
rect 1467 438 1535 472
rect 1625 438 1693 472
rect 1783 438 1851 472
rect 1941 438 2009 472
rect 2099 438 2167 472
rect 2257 438 2325 472
rect 2415 438 2483 472
rect 2573 438 2641 472
rect 2731 438 2799 472
rect 2889 438 2957 472
rect 3047 438 3115 472
rect 3205 438 3273 472
rect 3363 438 3431 472
rect 3521 438 3589 472
rect 3679 438 3747 472
rect 3837 438 3905 472
rect 3995 438 4063 472
rect 4153 438 4221 472
rect 4311 438 4379 472
rect 4469 438 4537 472
rect 4627 438 4695 472
rect 4785 438 4853 472
rect 4943 438 5011 472
rect 5101 438 5169 472
rect 5259 438 5327 472
rect 5417 438 5485 472
rect 5575 438 5643 472
rect 5733 438 5801 472
rect 5891 438 5959 472
rect 6049 438 6117 472
rect 6207 438 6275 472
rect -6275 -472 -6207 -438
rect -6117 -472 -6049 -438
rect -5959 -472 -5891 -438
rect -5801 -472 -5733 -438
rect -5643 -472 -5575 -438
rect -5485 -472 -5417 -438
rect -5327 -472 -5259 -438
rect -5169 -472 -5101 -438
rect -5011 -472 -4943 -438
rect -4853 -472 -4785 -438
rect -4695 -472 -4627 -438
rect -4537 -472 -4469 -438
rect -4379 -472 -4311 -438
rect -4221 -472 -4153 -438
rect -4063 -472 -3995 -438
rect -3905 -472 -3837 -438
rect -3747 -472 -3679 -438
rect -3589 -472 -3521 -438
rect -3431 -472 -3363 -438
rect -3273 -472 -3205 -438
rect -3115 -472 -3047 -438
rect -2957 -472 -2889 -438
rect -2799 -472 -2731 -438
rect -2641 -472 -2573 -438
rect -2483 -472 -2415 -438
rect -2325 -472 -2257 -438
rect -2167 -472 -2099 -438
rect -2009 -472 -1941 -438
rect -1851 -472 -1783 -438
rect -1693 -472 -1625 -438
rect -1535 -472 -1467 -438
rect -1377 -472 -1309 -438
rect -1219 -472 -1151 -438
rect -1061 -472 -993 -438
rect -903 -472 -835 -438
rect -745 -472 -677 -438
rect -587 -472 -519 -438
rect -429 -472 -361 -438
rect -271 -472 -203 -438
rect -113 -472 -45 -438
rect 45 -472 113 -438
rect 203 -472 271 -438
rect 361 -472 429 -438
rect 519 -472 587 -438
rect 677 -472 745 -438
rect 835 -472 903 -438
rect 993 -472 1061 -438
rect 1151 -472 1219 -438
rect 1309 -472 1377 -438
rect 1467 -472 1535 -438
rect 1625 -472 1693 -438
rect 1783 -472 1851 -438
rect 1941 -472 2009 -438
rect 2099 -472 2167 -438
rect 2257 -472 2325 -438
rect 2415 -472 2483 -438
rect 2573 -472 2641 -438
rect 2731 -472 2799 -438
rect 2889 -472 2957 -438
rect 3047 -472 3115 -438
rect 3205 -472 3273 -438
rect 3363 -472 3431 -438
rect 3521 -472 3589 -438
rect 3679 -472 3747 -438
rect 3837 -472 3905 -438
rect 3995 -472 4063 -438
rect 4153 -472 4221 -438
rect 4311 -472 4379 -438
rect 4469 -472 4537 -438
rect 4627 -472 4695 -438
rect 4785 -472 4853 -438
rect 4943 -472 5011 -438
rect 5101 -472 5169 -438
rect 5259 -472 5327 -438
rect 5417 -472 5485 -438
rect 5575 -472 5643 -438
rect 5733 -472 5801 -438
rect 5891 -472 5959 -438
rect 6049 -472 6117 -438
rect 6207 -472 6275 -438
<< locali >>
rect -6471 576 -6375 610
rect 6375 576 6471 610
rect -6471 514 -6437 576
rect 6437 514 6471 576
rect -6291 438 -6275 472
rect -6207 438 -6191 472
rect -6133 438 -6117 472
rect -6049 438 -6033 472
rect -5975 438 -5959 472
rect -5891 438 -5875 472
rect -5817 438 -5801 472
rect -5733 438 -5717 472
rect -5659 438 -5643 472
rect -5575 438 -5559 472
rect -5501 438 -5485 472
rect -5417 438 -5401 472
rect -5343 438 -5327 472
rect -5259 438 -5243 472
rect -5185 438 -5169 472
rect -5101 438 -5085 472
rect -5027 438 -5011 472
rect -4943 438 -4927 472
rect -4869 438 -4853 472
rect -4785 438 -4769 472
rect -4711 438 -4695 472
rect -4627 438 -4611 472
rect -4553 438 -4537 472
rect -4469 438 -4453 472
rect -4395 438 -4379 472
rect -4311 438 -4295 472
rect -4237 438 -4221 472
rect -4153 438 -4137 472
rect -4079 438 -4063 472
rect -3995 438 -3979 472
rect -3921 438 -3905 472
rect -3837 438 -3821 472
rect -3763 438 -3747 472
rect -3679 438 -3663 472
rect -3605 438 -3589 472
rect -3521 438 -3505 472
rect -3447 438 -3431 472
rect -3363 438 -3347 472
rect -3289 438 -3273 472
rect -3205 438 -3189 472
rect -3131 438 -3115 472
rect -3047 438 -3031 472
rect -2973 438 -2957 472
rect -2889 438 -2873 472
rect -2815 438 -2799 472
rect -2731 438 -2715 472
rect -2657 438 -2641 472
rect -2573 438 -2557 472
rect -2499 438 -2483 472
rect -2415 438 -2399 472
rect -2341 438 -2325 472
rect -2257 438 -2241 472
rect -2183 438 -2167 472
rect -2099 438 -2083 472
rect -2025 438 -2009 472
rect -1941 438 -1925 472
rect -1867 438 -1851 472
rect -1783 438 -1767 472
rect -1709 438 -1693 472
rect -1625 438 -1609 472
rect -1551 438 -1535 472
rect -1467 438 -1451 472
rect -1393 438 -1377 472
rect -1309 438 -1293 472
rect -1235 438 -1219 472
rect -1151 438 -1135 472
rect -1077 438 -1061 472
rect -993 438 -977 472
rect -919 438 -903 472
rect -835 438 -819 472
rect -761 438 -745 472
rect -677 438 -661 472
rect -603 438 -587 472
rect -519 438 -503 472
rect -445 438 -429 472
rect -361 438 -345 472
rect -287 438 -271 472
rect -203 438 -187 472
rect -129 438 -113 472
rect -45 438 -29 472
rect 29 438 45 472
rect 113 438 129 472
rect 187 438 203 472
rect 271 438 287 472
rect 345 438 361 472
rect 429 438 445 472
rect 503 438 519 472
rect 587 438 603 472
rect 661 438 677 472
rect 745 438 761 472
rect 819 438 835 472
rect 903 438 919 472
rect 977 438 993 472
rect 1061 438 1077 472
rect 1135 438 1151 472
rect 1219 438 1235 472
rect 1293 438 1309 472
rect 1377 438 1393 472
rect 1451 438 1467 472
rect 1535 438 1551 472
rect 1609 438 1625 472
rect 1693 438 1709 472
rect 1767 438 1783 472
rect 1851 438 1867 472
rect 1925 438 1941 472
rect 2009 438 2025 472
rect 2083 438 2099 472
rect 2167 438 2183 472
rect 2241 438 2257 472
rect 2325 438 2341 472
rect 2399 438 2415 472
rect 2483 438 2499 472
rect 2557 438 2573 472
rect 2641 438 2657 472
rect 2715 438 2731 472
rect 2799 438 2815 472
rect 2873 438 2889 472
rect 2957 438 2973 472
rect 3031 438 3047 472
rect 3115 438 3131 472
rect 3189 438 3205 472
rect 3273 438 3289 472
rect 3347 438 3363 472
rect 3431 438 3447 472
rect 3505 438 3521 472
rect 3589 438 3605 472
rect 3663 438 3679 472
rect 3747 438 3763 472
rect 3821 438 3837 472
rect 3905 438 3921 472
rect 3979 438 3995 472
rect 4063 438 4079 472
rect 4137 438 4153 472
rect 4221 438 4237 472
rect 4295 438 4311 472
rect 4379 438 4395 472
rect 4453 438 4469 472
rect 4537 438 4553 472
rect 4611 438 4627 472
rect 4695 438 4711 472
rect 4769 438 4785 472
rect 4853 438 4869 472
rect 4927 438 4943 472
rect 5011 438 5027 472
rect 5085 438 5101 472
rect 5169 438 5185 472
rect 5243 438 5259 472
rect 5327 438 5343 472
rect 5401 438 5417 472
rect 5485 438 5501 472
rect 5559 438 5575 472
rect 5643 438 5659 472
rect 5717 438 5733 472
rect 5801 438 5817 472
rect 5875 438 5891 472
rect 5959 438 5975 472
rect 6033 438 6049 472
rect 6117 438 6133 472
rect 6191 438 6207 472
rect 6275 438 6291 472
rect -6337 388 -6303 404
rect -6337 -404 -6303 -388
rect -6179 388 -6145 404
rect -6179 -404 -6145 -388
rect -6021 388 -5987 404
rect -6021 -404 -5987 -388
rect -5863 388 -5829 404
rect -5863 -404 -5829 -388
rect -5705 388 -5671 404
rect -5705 -404 -5671 -388
rect -5547 388 -5513 404
rect -5547 -404 -5513 -388
rect -5389 388 -5355 404
rect -5389 -404 -5355 -388
rect -5231 388 -5197 404
rect -5231 -404 -5197 -388
rect -5073 388 -5039 404
rect -5073 -404 -5039 -388
rect -4915 388 -4881 404
rect -4915 -404 -4881 -388
rect -4757 388 -4723 404
rect -4757 -404 -4723 -388
rect -4599 388 -4565 404
rect -4599 -404 -4565 -388
rect -4441 388 -4407 404
rect -4441 -404 -4407 -388
rect -4283 388 -4249 404
rect -4283 -404 -4249 -388
rect -4125 388 -4091 404
rect -4125 -404 -4091 -388
rect -3967 388 -3933 404
rect -3967 -404 -3933 -388
rect -3809 388 -3775 404
rect -3809 -404 -3775 -388
rect -3651 388 -3617 404
rect -3651 -404 -3617 -388
rect -3493 388 -3459 404
rect -3493 -404 -3459 -388
rect -3335 388 -3301 404
rect -3335 -404 -3301 -388
rect -3177 388 -3143 404
rect -3177 -404 -3143 -388
rect -3019 388 -2985 404
rect -3019 -404 -2985 -388
rect -2861 388 -2827 404
rect -2861 -404 -2827 -388
rect -2703 388 -2669 404
rect -2703 -404 -2669 -388
rect -2545 388 -2511 404
rect -2545 -404 -2511 -388
rect -2387 388 -2353 404
rect -2387 -404 -2353 -388
rect -2229 388 -2195 404
rect -2229 -404 -2195 -388
rect -2071 388 -2037 404
rect -2071 -404 -2037 -388
rect -1913 388 -1879 404
rect -1913 -404 -1879 -388
rect -1755 388 -1721 404
rect -1755 -404 -1721 -388
rect -1597 388 -1563 404
rect -1597 -404 -1563 -388
rect -1439 388 -1405 404
rect -1439 -404 -1405 -388
rect -1281 388 -1247 404
rect -1281 -404 -1247 -388
rect -1123 388 -1089 404
rect -1123 -404 -1089 -388
rect -965 388 -931 404
rect -965 -404 -931 -388
rect -807 388 -773 404
rect -807 -404 -773 -388
rect -649 388 -615 404
rect -649 -404 -615 -388
rect -491 388 -457 404
rect -491 -404 -457 -388
rect -333 388 -299 404
rect -333 -404 -299 -388
rect -175 388 -141 404
rect -175 -404 -141 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 141 388 175 404
rect 141 -404 175 -388
rect 299 388 333 404
rect 299 -404 333 -388
rect 457 388 491 404
rect 457 -404 491 -388
rect 615 388 649 404
rect 615 -404 649 -388
rect 773 388 807 404
rect 773 -404 807 -388
rect 931 388 965 404
rect 931 -404 965 -388
rect 1089 388 1123 404
rect 1089 -404 1123 -388
rect 1247 388 1281 404
rect 1247 -404 1281 -388
rect 1405 388 1439 404
rect 1405 -404 1439 -388
rect 1563 388 1597 404
rect 1563 -404 1597 -388
rect 1721 388 1755 404
rect 1721 -404 1755 -388
rect 1879 388 1913 404
rect 1879 -404 1913 -388
rect 2037 388 2071 404
rect 2037 -404 2071 -388
rect 2195 388 2229 404
rect 2195 -404 2229 -388
rect 2353 388 2387 404
rect 2353 -404 2387 -388
rect 2511 388 2545 404
rect 2511 -404 2545 -388
rect 2669 388 2703 404
rect 2669 -404 2703 -388
rect 2827 388 2861 404
rect 2827 -404 2861 -388
rect 2985 388 3019 404
rect 2985 -404 3019 -388
rect 3143 388 3177 404
rect 3143 -404 3177 -388
rect 3301 388 3335 404
rect 3301 -404 3335 -388
rect 3459 388 3493 404
rect 3459 -404 3493 -388
rect 3617 388 3651 404
rect 3617 -404 3651 -388
rect 3775 388 3809 404
rect 3775 -404 3809 -388
rect 3933 388 3967 404
rect 3933 -404 3967 -388
rect 4091 388 4125 404
rect 4091 -404 4125 -388
rect 4249 388 4283 404
rect 4249 -404 4283 -388
rect 4407 388 4441 404
rect 4407 -404 4441 -388
rect 4565 388 4599 404
rect 4565 -404 4599 -388
rect 4723 388 4757 404
rect 4723 -404 4757 -388
rect 4881 388 4915 404
rect 4881 -404 4915 -388
rect 5039 388 5073 404
rect 5039 -404 5073 -388
rect 5197 388 5231 404
rect 5197 -404 5231 -388
rect 5355 388 5389 404
rect 5355 -404 5389 -388
rect 5513 388 5547 404
rect 5513 -404 5547 -388
rect 5671 388 5705 404
rect 5671 -404 5705 -388
rect 5829 388 5863 404
rect 5829 -404 5863 -388
rect 5987 388 6021 404
rect 5987 -404 6021 -388
rect 6145 388 6179 404
rect 6145 -404 6179 -388
rect 6303 388 6337 404
rect 6303 -404 6337 -388
rect -6291 -472 -6275 -438
rect -6207 -472 -6191 -438
rect -6133 -472 -6117 -438
rect -6049 -472 -6033 -438
rect -5975 -472 -5959 -438
rect -5891 -472 -5875 -438
rect -5817 -472 -5801 -438
rect -5733 -472 -5717 -438
rect -5659 -472 -5643 -438
rect -5575 -472 -5559 -438
rect -5501 -472 -5485 -438
rect -5417 -472 -5401 -438
rect -5343 -472 -5327 -438
rect -5259 -472 -5243 -438
rect -5185 -472 -5169 -438
rect -5101 -472 -5085 -438
rect -5027 -472 -5011 -438
rect -4943 -472 -4927 -438
rect -4869 -472 -4853 -438
rect -4785 -472 -4769 -438
rect -4711 -472 -4695 -438
rect -4627 -472 -4611 -438
rect -4553 -472 -4537 -438
rect -4469 -472 -4453 -438
rect -4395 -472 -4379 -438
rect -4311 -472 -4295 -438
rect -4237 -472 -4221 -438
rect -4153 -472 -4137 -438
rect -4079 -472 -4063 -438
rect -3995 -472 -3979 -438
rect -3921 -472 -3905 -438
rect -3837 -472 -3821 -438
rect -3763 -472 -3747 -438
rect -3679 -472 -3663 -438
rect -3605 -472 -3589 -438
rect -3521 -472 -3505 -438
rect -3447 -472 -3431 -438
rect -3363 -472 -3347 -438
rect -3289 -472 -3273 -438
rect -3205 -472 -3189 -438
rect -3131 -472 -3115 -438
rect -3047 -472 -3031 -438
rect -2973 -472 -2957 -438
rect -2889 -472 -2873 -438
rect -2815 -472 -2799 -438
rect -2731 -472 -2715 -438
rect -2657 -472 -2641 -438
rect -2573 -472 -2557 -438
rect -2499 -472 -2483 -438
rect -2415 -472 -2399 -438
rect -2341 -472 -2325 -438
rect -2257 -472 -2241 -438
rect -2183 -472 -2167 -438
rect -2099 -472 -2083 -438
rect -2025 -472 -2009 -438
rect -1941 -472 -1925 -438
rect -1867 -472 -1851 -438
rect -1783 -472 -1767 -438
rect -1709 -472 -1693 -438
rect -1625 -472 -1609 -438
rect -1551 -472 -1535 -438
rect -1467 -472 -1451 -438
rect -1393 -472 -1377 -438
rect -1309 -472 -1293 -438
rect -1235 -472 -1219 -438
rect -1151 -472 -1135 -438
rect -1077 -472 -1061 -438
rect -993 -472 -977 -438
rect -919 -472 -903 -438
rect -835 -472 -819 -438
rect -761 -472 -745 -438
rect -677 -472 -661 -438
rect -603 -472 -587 -438
rect -519 -472 -503 -438
rect -445 -472 -429 -438
rect -361 -472 -345 -438
rect -287 -472 -271 -438
rect -203 -472 -187 -438
rect -129 -472 -113 -438
rect -45 -472 -29 -438
rect 29 -472 45 -438
rect 113 -472 129 -438
rect 187 -472 203 -438
rect 271 -472 287 -438
rect 345 -472 361 -438
rect 429 -472 445 -438
rect 503 -472 519 -438
rect 587 -472 603 -438
rect 661 -472 677 -438
rect 745 -472 761 -438
rect 819 -472 835 -438
rect 903 -472 919 -438
rect 977 -472 993 -438
rect 1061 -472 1077 -438
rect 1135 -472 1151 -438
rect 1219 -472 1235 -438
rect 1293 -472 1309 -438
rect 1377 -472 1393 -438
rect 1451 -472 1467 -438
rect 1535 -472 1551 -438
rect 1609 -472 1625 -438
rect 1693 -472 1709 -438
rect 1767 -472 1783 -438
rect 1851 -472 1867 -438
rect 1925 -472 1941 -438
rect 2009 -472 2025 -438
rect 2083 -472 2099 -438
rect 2167 -472 2183 -438
rect 2241 -472 2257 -438
rect 2325 -472 2341 -438
rect 2399 -472 2415 -438
rect 2483 -472 2499 -438
rect 2557 -472 2573 -438
rect 2641 -472 2657 -438
rect 2715 -472 2731 -438
rect 2799 -472 2815 -438
rect 2873 -472 2889 -438
rect 2957 -472 2973 -438
rect 3031 -472 3047 -438
rect 3115 -472 3131 -438
rect 3189 -472 3205 -438
rect 3273 -472 3289 -438
rect 3347 -472 3363 -438
rect 3431 -472 3447 -438
rect 3505 -472 3521 -438
rect 3589 -472 3605 -438
rect 3663 -472 3679 -438
rect 3747 -472 3763 -438
rect 3821 -472 3837 -438
rect 3905 -472 3921 -438
rect 3979 -472 3995 -438
rect 4063 -472 4079 -438
rect 4137 -472 4153 -438
rect 4221 -472 4237 -438
rect 4295 -472 4311 -438
rect 4379 -472 4395 -438
rect 4453 -472 4469 -438
rect 4537 -472 4553 -438
rect 4611 -472 4627 -438
rect 4695 -472 4711 -438
rect 4769 -472 4785 -438
rect 4853 -472 4869 -438
rect 4927 -472 4943 -438
rect 5011 -472 5027 -438
rect 5085 -472 5101 -438
rect 5169 -472 5185 -438
rect 5243 -472 5259 -438
rect 5327 -472 5343 -438
rect 5401 -472 5417 -438
rect 5485 -472 5501 -438
rect 5559 -472 5575 -438
rect 5643 -472 5659 -438
rect 5717 -472 5733 -438
rect 5801 -472 5817 -438
rect 5875 -472 5891 -438
rect 5959 -472 5975 -438
rect 6033 -472 6049 -438
rect 6117 -472 6133 -438
rect 6191 -472 6207 -438
rect 6275 -472 6291 -438
rect -6471 -576 -6437 -514
rect 6437 -576 6471 -514
rect -6471 -610 -6375 -576
rect 6375 -610 6471 -576
<< viali >>
rect -6275 438 -6207 472
rect -6117 438 -6049 472
rect -5959 438 -5891 472
rect -5801 438 -5733 472
rect -5643 438 -5575 472
rect -5485 438 -5417 472
rect -5327 438 -5259 472
rect -5169 438 -5101 472
rect -5011 438 -4943 472
rect -4853 438 -4785 472
rect -4695 438 -4627 472
rect -4537 438 -4469 472
rect -4379 438 -4311 472
rect -4221 438 -4153 472
rect -4063 438 -3995 472
rect -3905 438 -3837 472
rect -3747 438 -3679 472
rect -3589 438 -3521 472
rect -3431 438 -3363 472
rect -3273 438 -3205 472
rect -3115 438 -3047 472
rect -2957 438 -2889 472
rect -2799 438 -2731 472
rect -2641 438 -2573 472
rect -2483 438 -2415 472
rect -2325 438 -2257 472
rect -2167 438 -2099 472
rect -2009 438 -1941 472
rect -1851 438 -1783 472
rect -1693 438 -1625 472
rect -1535 438 -1467 472
rect -1377 438 -1309 472
rect -1219 438 -1151 472
rect -1061 438 -993 472
rect -903 438 -835 472
rect -745 438 -677 472
rect -587 438 -519 472
rect -429 438 -361 472
rect -271 438 -203 472
rect -113 438 -45 472
rect 45 438 113 472
rect 203 438 271 472
rect 361 438 429 472
rect 519 438 587 472
rect 677 438 745 472
rect 835 438 903 472
rect 993 438 1061 472
rect 1151 438 1219 472
rect 1309 438 1377 472
rect 1467 438 1535 472
rect 1625 438 1693 472
rect 1783 438 1851 472
rect 1941 438 2009 472
rect 2099 438 2167 472
rect 2257 438 2325 472
rect 2415 438 2483 472
rect 2573 438 2641 472
rect 2731 438 2799 472
rect 2889 438 2957 472
rect 3047 438 3115 472
rect 3205 438 3273 472
rect 3363 438 3431 472
rect 3521 438 3589 472
rect 3679 438 3747 472
rect 3837 438 3905 472
rect 3995 438 4063 472
rect 4153 438 4221 472
rect 4311 438 4379 472
rect 4469 438 4537 472
rect 4627 438 4695 472
rect 4785 438 4853 472
rect 4943 438 5011 472
rect 5101 438 5169 472
rect 5259 438 5327 472
rect 5417 438 5485 472
rect 5575 438 5643 472
rect 5733 438 5801 472
rect 5891 438 5959 472
rect 6049 438 6117 472
rect 6207 438 6275 472
rect -6337 -388 -6303 388
rect -6179 -388 -6145 388
rect -6021 -388 -5987 388
rect -5863 -388 -5829 388
rect -5705 -388 -5671 388
rect -5547 -388 -5513 388
rect -5389 -388 -5355 388
rect -5231 -388 -5197 388
rect -5073 -388 -5039 388
rect -4915 -388 -4881 388
rect -4757 -388 -4723 388
rect -4599 -388 -4565 388
rect -4441 -388 -4407 388
rect -4283 -388 -4249 388
rect -4125 -388 -4091 388
rect -3967 -388 -3933 388
rect -3809 -388 -3775 388
rect -3651 -388 -3617 388
rect -3493 -388 -3459 388
rect -3335 -388 -3301 388
rect -3177 -388 -3143 388
rect -3019 -388 -2985 388
rect -2861 -388 -2827 388
rect -2703 -388 -2669 388
rect -2545 -388 -2511 388
rect -2387 -388 -2353 388
rect -2229 -388 -2195 388
rect -2071 -388 -2037 388
rect -1913 -388 -1879 388
rect -1755 -388 -1721 388
rect -1597 -388 -1563 388
rect -1439 -388 -1405 388
rect -1281 -388 -1247 388
rect -1123 -388 -1089 388
rect -965 -388 -931 388
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
rect 931 -388 965 388
rect 1089 -388 1123 388
rect 1247 -388 1281 388
rect 1405 -388 1439 388
rect 1563 -388 1597 388
rect 1721 -388 1755 388
rect 1879 -388 1913 388
rect 2037 -388 2071 388
rect 2195 -388 2229 388
rect 2353 -388 2387 388
rect 2511 -388 2545 388
rect 2669 -388 2703 388
rect 2827 -388 2861 388
rect 2985 -388 3019 388
rect 3143 -388 3177 388
rect 3301 -388 3335 388
rect 3459 -388 3493 388
rect 3617 -388 3651 388
rect 3775 -388 3809 388
rect 3933 -388 3967 388
rect 4091 -388 4125 388
rect 4249 -388 4283 388
rect 4407 -388 4441 388
rect 4565 -388 4599 388
rect 4723 -388 4757 388
rect 4881 -388 4915 388
rect 5039 -388 5073 388
rect 5197 -388 5231 388
rect 5355 -388 5389 388
rect 5513 -388 5547 388
rect 5671 -388 5705 388
rect 5829 -388 5863 388
rect 5987 -388 6021 388
rect 6145 -388 6179 388
rect 6303 -388 6337 388
rect -6275 -472 -6207 -438
rect -6117 -472 -6049 -438
rect -5959 -472 -5891 -438
rect -5801 -472 -5733 -438
rect -5643 -472 -5575 -438
rect -5485 -472 -5417 -438
rect -5327 -472 -5259 -438
rect -5169 -472 -5101 -438
rect -5011 -472 -4943 -438
rect -4853 -472 -4785 -438
rect -4695 -472 -4627 -438
rect -4537 -472 -4469 -438
rect -4379 -472 -4311 -438
rect -4221 -472 -4153 -438
rect -4063 -472 -3995 -438
rect -3905 -472 -3837 -438
rect -3747 -472 -3679 -438
rect -3589 -472 -3521 -438
rect -3431 -472 -3363 -438
rect -3273 -472 -3205 -438
rect -3115 -472 -3047 -438
rect -2957 -472 -2889 -438
rect -2799 -472 -2731 -438
rect -2641 -472 -2573 -438
rect -2483 -472 -2415 -438
rect -2325 -472 -2257 -438
rect -2167 -472 -2099 -438
rect -2009 -472 -1941 -438
rect -1851 -472 -1783 -438
rect -1693 -472 -1625 -438
rect -1535 -472 -1467 -438
rect -1377 -472 -1309 -438
rect -1219 -472 -1151 -438
rect -1061 -472 -993 -438
rect -903 -472 -835 -438
rect -745 -472 -677 -438
rect -587 -472 -519 -438
rect -429 -472 -361 -438
rect -271 -472 -203 -438
rect -113 -472 -45 -438
rect 45 -472 113 -438
rect 203 -472 271 -438
rect 361 -472 429 -438
rect 519 -472 587 -438
rect 677 -472 745 -438
rect 835 -472 903 -438
rect 993 -472 1061 -438
rect 1151 -472 1219 -438
rect 1309 -472 1377 -438
rect 1467 -472 1535 -438
rect 1625 -472 1693 -438
rect 1783 -472 1851 -438
rect 1941 -472 2009 -438
rect 2099 -472 2167 -438
rect 2257 -472 2325 -438
rect 2415 -472 2483 -438
rect 2573 -472 2641 -438
rect 2731 -472 2799 -438
rect 2889 -472 2957 -438
rect 3047 -472 3115 -438
rect 3205 -472 3273 -438
rect 3363 -472 3431 -438
rect 3521 -472 3589 -438
rect 3679 -472 3747 -438
rect 3837 -472 3905 -438
rect 3995 -472 4063 -438
rect 4153 -472 4221 -438
rect 4311 -472 4379 -438
rect 4469 -472 4537 -438
rect 4627 -472 4695 -438
rect 4785 -472 4853 -438
rect 4943 -472 5011 -438
rect 5101 -472 5169 -438
rect 5259 -472 5327 -438
rect 5417 -472 5485 -438
rect 5575 -472 5643 -438
rect 5733 -472 5801 -438
rect 5891 -472 5959 -438
rect 6049 -472 6117 -438
rect 6207 -472 6275 -438
<< metal1 >>
rect -6287 472 -6195 478
rect -6287 438 -6275 472
rect -6207 438 -6195 472
rect -6287 432 -6195 438
rect -6129 472 -6037 478
rect -6129 438 -6117 472
rect -6049 438 -6037 472
rect -6129 432 -6037 438
rect -5971 472 -5879 478
rect -5971 438 -5959 472
rect -5891 438 -5879 472
rect -5971 432 -5879 438
rect -5813 472 -5721 478
rect -5813 438 -5801 472
rect -5733 438 -5721 472
rect -5813 432 -5721 438
rect -5655 472 -5563 478
rect -5655 438 -5643 472
rect -5575 438 -5563 472
rect -5655 432 -5563 438
rect -5497 472 -5405 478
rect -5497 438 -5485 472
rect -5417 438 -5405 472
rect -5497 432 -5405 438
rect -5339 472 -5247 478
rect -5339 438 -5327 472
rect -5259 438 -5247 472
rect -5339 432 -5247 438
rect -5181 472 -5089 478
rect -5181 438 -5169 472
rect -5101 438 -5089 472
rect -5181 432 -5089 438
rect -5023 472 -4931 478
rect -5023 438 -5011 472
rect -4943 438 -4931 472
rect -5023 432 -4931 438
rect -4865 472 -4773 478
rect -4865 438 -4853 472
rect -4785 438 -4773 472
rect -4865 432 -4773 438
rect -4707 472 -4615 478
rect -4707 438 -4695 472
rect -4627 438 -4615 472
rect -4707 432 -4615 438
rect -4549 472 -4457 478
rect -4549 438 -4537 472
rect -4469 438 -4457 472
rect -4549 432 -4457 438
rect -4391 472 -4299 478
rect -4391 438 -4379 472
rect -4311 438 -4299 472
rect -4391 432 -4299 438
rect -4233 472 -4141 478
rect -4233 438 -4221 472
rect -4153 438 -4141 472
rect -4233 432 -4141 438
rect -4075 472 -3983 478
rect -4075 438 -4063 472
rect -3995 438 -3983 472
rect -4075 432 -3983 438
rect -3917 472 -3825 478
rect -3917 438 -3905 472
rect -3837 438 -3825 472
rect -3917 432 -3825 438
rect -3759 472 -3667 478
rect -3759 438 -3747 472
rect -3679 438 -3667 472
rect -3759 432 -3667 438
rect -3601 472 -3509 478
rect -3601 438 -3589 472
rect -3521 438 -3509 472
rect -3601 432 -3509 438
rect -3443 472 -3351 478
rect -3443 438 -3431 472
rect -3363 438 -3351 472
rect -3443 432 -3351 438
rect -3285 472 -3193 478
rect -3285 438 -3273 472
rect -3205 438 -3193 472
rect -3285 432 -3193 438
rect -3127 472 -3035 478
rect -3127 438 -3115 472
rect -3047 438 -3035 472
rect -3127 432 -3035 438
rect -2969 472 -2877 478
rect -2969 438 -2957 472
rect -2889 438 -2877 472
rect -2969 432 -2877 438
rect -2811 472 -2719 478
rect -2811 438 -2799 472
rect -2731 438 -2719 472
rect -2811 432 -2719 438
rect -2653 472 -2561 478
rect -2653 438 -2641 472
rect -2573 438 -2561 472
rect -2653 432 -2561 438
rect -2495 472 -2403 478
rect -2495 438 -2483 472
rect -2415 438 -2403 472
rect -2495 432 -2403 438
rect -2337 472 -2245 478
rect -2337 438 -2325 472
rect -2257 438 -2245 472
rect -2337 432 -2245 438
rect -2179 472 -2087 478
rect -2179 438 -2167 472
rect -2099 438 -2087 472
rect -2179 432 -2087 438
rect -2021 472 -1929 478
rect -2021 438 -2009 472
rect -1941 438 -1929 472
rect -2021 432 -1929 438
rect -1863 472 -1771 478
rect -1863 438 -1851 472
rect -1783 438 -1771 472
rect -1863 432 -1771 438
rect -1705 472 -1613 478
rect -1705 438 -1693 472
rect -1625 438 -1613 472
rect -1705 432 -1613 438
rect -1547 472 -1455 478
rect -1547 438 -1535 472
rect -1467 438 -1455 472
rect -1547 432 -1455 438
rect -1389 472 -1297 478
rect -1389 438 -1377 472
rect -1309 438 -1297 472
rect -1389 432 -1297 438
rect -1231 472 -1139 478
rect -1231 438 -1219 472
rect -1151 438 -1139 472
rect -1231 432 -1139 438
rect -1073 472 -981 478
rect -1073 438 -1061 472
rect -993 438 -981 472
rect -1073 432 -981 438
rect -915 472 -823 478
rect -915 438 -903 472
rect -835 438 -823 472
rect -915 432 -823 438
rect -757 472 -665 478
rect -757 438 -745 472
rect -677 438 -665 472
rect -757 432 -665 438
rect -599 472 -507 478
rect -599 438 -587 472
rect -519 438 -507 472
rect -599 432 -507 438
rect -441 472 -349 478
rect -441 438 -429 472
rect -361 438 -349 472
rect -441 432 -349 438
rect -283 472 -191 478
rect -283 438 -271 472
rect -203 438 -191 472
rect -283 432 -191 438
rect -125 472 -33 478
rect -125 438 -113 472
rect -45 438 -33 472
rect -125 432 -33 438
rect 33 472 125 478
rect 33 438 45 472
rect 113 438 125 472
rect 33 432 125 438
rect 191 472 283 478
rect 191 438 203 472
rect 271 438 283 472
rect 191 432 283 438
rect 349 472 441 478
rect 349 438 361 472
rect 429 438 441 472
rect 349 432 441 438
rect 507 472 599 478
rect 507 438 519 472
rect 587 438 599 472
rect 507 432 599 438
rect 665 472 757 478
rect 665 438 677 472
rect 745 438 757 472
rect 665 432 757 438
rect 823 472 915 478
rect 823 438 835 472
rect 903 438 915 472
rect 823 432 915 438
rect 981 472 1073 478
rect 981 438 993 472
rect 1061 438 1073 472
rect 981 432 1073 438
rect 1139 472 1231 478
rect 1139 438 1151 472
rect 1219 438 1231 472
rect 1139 432 1231 438
rect 1297 472 1389 478
rect 1297 438 1309 472
rect 1377 438 1389 472
rect 1297 432 1389 438
rect 1455 472 1547 478
rect 1455 438 1467 472
rect 1535 438 1547 472
rect 1455 432 1547 438
rect 1613 472 1705 478
rect 1613 438 1625 472
rect 1693 438 1705 472
rect 1613 432 1705 438
rect 1771 472 1863 478
rect 1771 438 1783 472
rect 1851 438 1863 472
rect 1771 432 1863 438
rect 1929 472 2021 478
rect 1929 438 1941 472
rect 2009 438 2021 472
rect 1929 432 2021 438
rect 2087 472 2179 478
rect 2087 438 2099 472
rect 2167 438 2179 472
rect 2087 432 2179 438
rect 2245 472 2337 478
rect 2245 438 2257 472
rect 2325 438 2337 472
rect 2245 432 2337 438
rect 2403 472 2495 478
rect 2403 438 2415 472
rect 2483 438 2495 472
rect 2403 432 2495 438
rect 2561 472 2653 478
rect 2561 438 2573 472
rect 2641 438 2653 472
rect 2561 432 2653 438
rect 2719 472 2811 478
rect 2719 438 2731 472
rect 2799 438 2811 472
rect 2719 432 2811 438
rect 2877 472 2969 478
rect 2877 438 2889 472
rect 2957 438 2969 472
rect 2877 432 2969 438
rect 3035 472 3127 478
rect 3035 438 3047 472
rect 3115 438 3127 472
rect 3035 432 3127 438
rect 3193 472 3285 478
rect 3193 438 3205 472
rect 3273 438 3285 472
rect 3193 432 3285 438
rect 3351 472 3443 478
rect 3351 438 3363 472
rect 3431 438 3443 472
rect 3351 432 3443 438
rect 3509 472 3601 478
rect 3509 438 3521 472
rect 3589 438 3601 472
rect 3509 432 3601 438
rect 3667 472 3759 478
rect 3667 438 3679 472
rect 3747 438 3759 472
rect 3667 432 3759 438
rect 3825 472 3917 478
rect 3825 438 3837 472
rect 3905 438 3917 472
rect 3825 432 3917 438
rect 3983 472 4075 478
rect 3983 438 3995 472
rect 4063 438 4075 472
rect 3983 432 4075 438
rect 4141 472 4233 478
rect 4141 438 4153 472
rect 4221 438 4233 472
rect 4141 432 4233 438
rect 4299 472 4391 478
rect 4299 438 4311 472
rect 4379 438 4391 472
rect 4299 432 4391 438
rect 4457 472 4549 478
rect 4457 438 4469 472
rect 4537 438 4549 472
rect 4457 432 4549 438
rect 4615 472 4707 478
rect 4615 438 4627 472
rect 4695 438 4707 472
rect 4615 432 4707 438
rect 4773 472 4865 478
rect 4773 438 4785 472
rect 4853 438 4865 472
rect 4773 432 4865 438
rect 4931 472 5023 478
rect 4931 438 4943 472
rect 5011 438 5023 472
rect 4931 432 5023 438
rect 5089 472 5181 478
rect 5089 438 5101 472
rect 5169 438 5181 472
rect 5089 432 5181 438
rect 5247 472 5339 478
rect 5247 438 5259 472
rect 5327 438 5339 472
rect 5247 432 5339 438
rect 5405 472 5497 478
rect 5405 438 5417 472
rect 5485 438 5497 472
rect 5405 432 5497 438
rect 5563 472 5655 478
rect 5563 438 5575 472
rect 5643 438 5655 472
rect 5563 432 5655 438
rect 5721 472 5813 478
rect 5721 438 5733 472
rect 5801 438 5813 472
rect 5721 432 5813 438
rect 5879 472 5971 478
rect 5879 438 5891 472
rect 5959 438 5971 472
rect 5879 432 5971 438
rect 6037 472 6129 478
rect 6037 438 6049 472
rect 6117 438 6129 472
rect 6037 432 6129 438
rect 6195 472 6287 478
rect 6195 438 6207 472
rect 6275 438 6287 472
rect 6195 432 6287 438
rect -6343 388 -6297 400
rect -6343 -388 -6337 388
rect -6303 -388 -6297 388
rect -6343 -400 -6297 -388
rect -6185 388 -6139 400
rect -6185 -388 -6179 388
rect -6145 -388 -6139 388
rect -6185 -400 -6139 -388
rect -6027 388 -5981 400
rect -6027 -388 -6021 388
rect -5987 -388 -5981 388
rect -6027 -400 -5981 -388
rect -5869 388 -5823 400
rect -5869 -388 -5863 388
rect -5829 -388 -5823 388
rect -5869 -400 -5823 -388
rect -5711 388 -5665 400
rect -5711 -388 -5705 388
rect -5671 -388 -5665 388
rect -5711 -400 -5665 -388
rect -5553 388 -5507 400
rect -5553 -388 -5547 388
rect -5513 -388 -5507 388
rect -5553 -400 -5507 -388
rect -5395 388 -5349 400
rect -5395 -388 -5389 388
rect -5355 -388 -5349 388
rect -5395 -400 -5349 -388
rect -5237 388 -5191 400
rect -5237 -388 -5231 388
rect -5197 -388 -5191 388
rect -5237 -400 -5191 -388
rect -5079 388 -5033 400
rect -5079 -388 -5073 388
rect -5039 -388 -5033 388
rect -5079 -400 -5033 -388
rect -4921 388 -4875 400
rect -4921 -388 -4915 388
rect -4881 -388 -4875 388
rect -4921 -400 -4875 -388
rect -4763 388 -4717 400
rect -4763 -388 -4757 388
rect -4723 -388 -4717 388
rect -4763 -400 -4717 -388
rect -4605 388 -4559 400
rect -4605 -388 -4599 388
rect -4565 -388 -4559 388
rect -4605 -400 -4559 -388
rect -4447 388 -4401 400
rect -4447 -388 -4441 388
rect -4407 -388 -4401 388
rect -4447 -400 -4401 -388
rect -4289 388 -4243 400
rect -4289 -388 -4283 388
rect -4249 -388 -4243 388
rect -4289 -400 -4243 -388
rect -4131 388 -4085 400
rect -4131 -388 -4125 388
rect -4091 -388 -4085 388
rect -4131 -400 -4085 -388
rect -3973 388 -3927 400
rect -3973 -388 -3967 388
rect -3933 -388 -3927 388
rect -3973 -400 -3927 -388
rect -3815 388 -3769 400
rect -3815 -388 -3809 388
rect -3775 -388 -3769 388
rect -3815 -400 -3769 -388
rect -3657 388 -3611 400
rect -3657 -388 -3651 388
rect -3617 -388 -3611 388
rect -3657 -400 -3611 -388
rect -3499 388 -3453 400
rect -3499 -388 -3493 388
rect -3459 -388 -3453 388
rect -3499 -400 -3453 -388
rect -3341 388 -3295 400
rect -3341 -388 -3335 388
rect -3301 -388 -3295 388
rect -3341 -400 -3295 -388
rect -3183 388 -3137 400
rect -3183 -388 -3177 388
rect -3143 -388 -3137 388
rect -3183 -400 -3137 -388
rect -3025 388 -2979 400
rect -3025 -388 -3019 388
rect -2985 -388 -2979 388
rect -3025 -400 -2979 -388
rect -2867 388 -2821 400
rect -2867 -388 -2861 388
rect -2827 -388 -2821 388
rect -2867 -400 -2821 -388
rect -2709 388 -2663 400
rect -2709 -388 -2703 388
rect -2669 -388 -2663 388
rect -2709 -400 -2663 -388
rect -2551 388 -2505 400
rect -2551 -388 -2545 388
rect -2511 -388 -2505 388
rect -2551 -400 -2505 -388
rect -2393 388 -2347 400
rect -2393 -388 -2387 388
rect -2353 -388 -2347 388
rect -2393 -400 -2347 -388
rect -2235 388 -2189 400
rect -2235 -388 -2229 388
rect -2195 -388 -2189 388
rect -2235 -400 -2189 -388
rect -2077 388 -2031 400
rect -2077 -388 -2071 388
rect -2037 -388 -2031 388
rect -2077 -400 -2031 -388
rect -1919 388 -1873 400
rect -1919 -388 -1913 388
rect -1879 -388 -1873 388
rect -1919 -400 -1873 -388
rect -1761 388 -1715 400
rect -1761 -388 -1755 388
rect -1721 -388 -1715 388
rect -1761 -400 -1715 -388
rect -1603 388 -1557 400
rect -1603 -388 -1597 388
rect -1563 -388 -1557 388
rect -1603 -400 -1557 -388
rect -1445 388 -1399 400
rect -1445 -388 -1439 388
rect -1405 -388 -1399 388
rect -1445 -400 -1399 -388
rect -1287 388 -1241 400
rect -1287 -388 -1281 388
rect -1247 -388 -1241 388
rect -1287 -400 -1241 -388
rect -1129 388 -1083 400
rect -1129 -388 -1123 388
rect -1089 -388 -1083 388
rect -1129 -400 -1083 -388
rect -971 388 -925 400
rect -971 -388 -965 388
rect -931 -388 -925 388
rect -971 -400 -925 -388
rect -813 388 -767 400
rect -813 -388 -807 388
rect -773 -388 -767 388
rect -813 -400 -767 -388
rect -655 388 -609 400
rect -655 -388 -649 388
rect -615 -388 -609 388
rect -655 -400 -609 -388
rect -497 388 -451 400
rect -497 -388 -491 388
rect -457 -388 -451 388
rect -497 -400 -451 -388
rect -339 388 -293 400
rect -339 -388 -333 388
rect -299 -388 -293 388
rect -339 -400 -293 -388
rect -181 388 -135 400
rect -181 -388 -175 388
rect -141 -388 -135 388
rect -181 -400 -135 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 135 388 181 400
rect 135 -388 141 388
rect 175 -388 181 388
rect 135 -400 181 -388
rect 293 388 339 400
rect 293 -388 299 388
rect 333 -388 339 388
rect 293 -400 339 -388
rect 451 388 497 400
rect 451 -388 457 388
rect 491 -388 497 388
rect 451 -400 497 -388
rect 609 388 655 400
rect 609 -388 615 388
rect 649 -388 655 388
rect 609 -400 655 -388
rect 767 388 813 400
rect 767 -388 773 388
rect 807 -388 813 388
rect 767 -400 813 -388
rect 925 388 971 400
rect 925 -388 931 388
rect 965 -388 971 388
rect 925 -400 971 -388
rect 1083 388 1129 400
rect 1083 -388 1089 388
rect 1123 -388 1129 388
rect 1083 -400 1129 -388
rect 1241 388 1287 400
rect 1241 -388 1247 388
rect 1281 -388 1287 388
rect 1241 -400 1287 -388
rect 1399 388 1445 400
rect 1399 -388 1405 388
rect 1439 -388 1445 388
rect 1399 -400 1445 -388
rect 1557 388 1603 400
rect 1557 -388 1563 388
rect 1597 -388 1603 388
rect 1557 -400 1603 -388
rect 1715 388 1761 400
rect 1715 -388 1721 388
rect 1755 -388 1761 388
rect 1715 -400 1761 -388
rect 1873 388 1919 400
rect 1873 -388 1879 388
rect 1913 -388 1919 388
rect 1873 -400 1919 -388
rect 2031 388 2077 400
rect 2031 -388 2037 388
rect 2071 -388 2077 388
rect 2031 -400 2077 -388
rect 2189 388 2235 400
rect 2189 -388 2195 388
rect 2229 -388 2235 388
rect 2189 -400 2235 -388
rect 2347 388 2393 400
rect 2347 -388 2353 388
rect 2387 -388 2393 388
rect 2347 -400 2393 -388
rect 2505 388 2551 400
rect 2505 -388 2511 388
rect 2545 -388 2551 388
rect 2505 -400 2551 -388
rect 2663 388 2709 400
rect 2663 -388 2669 388
rect 2703 -388 2709 388
rect 2663 -400 2709 -388
rect 2821 388 2867 400
rect 2821 -388 2827 388
rect 2861 -388 2867 388
rect 2821 -400 2867 -388
rect 2979 388 3025 400
rect 2979 -388 2985 388
rect 3019 -388 3025 388
rect 2979 -400 3025 -388
rect 3137 388 3183 400
rect 3137 -388 3143 388
rect 3177 -388 3183 388
rect 3137 -400 3183 -388
rect 3295 388 3341 400
rect 3295 -388 3301 388
rect 3335 -388 3341 388
rect 3295 -400 3341 -388
rect 3453 388 3499 400
rect 3453 -388 3459 388
rect 3493 -388 3499 388
rect 3453 -400 3499 -388
rect 3611 388 3657 400
rect 3611 -388 3617 388
rect 3651 -388 3657 388
rect 3611 -400 3657 -388
rect 3769 388 3815 400
rect 3769 -388 3775 388
rect 3809 -388 3815 388
rect 3769 -400 3815 -388
rect 3927 388 3973 400
rect 3927 -388 3933 388
rect 3967 -388 3973 388
rect 3927 -400 3973 -388
rect 4085 388 4131 400
rect 4085 -388 4091 388
rect 4125 -388 4131 388
rect 4085 -400 4131 -388
rect 4243 388 4289 400
rect 4243 -388 4249 388
rect 4283 -388 4289 388
rect 4243 -400 4289 -388
rect 4401 388 4447 400
rect 4401 -388 4407 388
rect 4441 -388 4447 388
rect 4401 -400 4447 -388
rect 4559 388 4605 400
rect 4559 -388 4565 388
rect 4599 -388 4605 388
rect 4559 -400 4605 -388
rect 4717 388 4763 400
rect 4717 -388 4723 388
rect 4757 -388 4763 388
rect 4717 -400 4763 -388
rect 4875 388 4921 400
rect 4875 -388 4881 388
rect 4915 -388 4921 388
rect 4875 -400 4921 -388
rect 5033 388 5079 400
rect 5033 -388 5039 388
rect 5073 -388 5079 388
rect 5033 -400 5079 -388
rect 5191 388 5237 400
rect 5191 -388 5197 388
rect 5231 -388 5237 388
rect 5191 -400 5237 -388
rect 5349 388 5395 400
rect 5349 -388 5355 388
rect 5389 -388 5395 388
rect 5349 -400 5395 -388
rect 5507 388 5553 400
rect 5507 -388 5513 388
rect 5547 -388 5553 388
rect 5507 -400 5553 -388
rect 5665 388 5711 400
rect 5665 -388 5671 388
rect 5705 -388 5711 388
rect 5665 -400 5711 -388
rect 5823 388 5869 400
rect 5823 -388 5829 388
rect 5863 -388 5869 388
rect 5823 -400 5869 -388
rect 5981 388 6027 400
rect 5981 -388 5987 388
rect 6021 -388 6027 388
rect 5981 -400 6027 -388
rect 6139 388 6185 400
rect 6139 -388 6145 388
rect 6179 -388 6185 388
rect 6139 -400 6185 -388
rect 6297 388 6343 400
rect 6297 -388 6303 388
rect 6337 -388 6343 388
rect 6297 -400 6343 -388
rect -6287 -438 -6195 -432
rect -6287 -472 -6275 -438
rect -6207 -472 -6195 -438
rect -6287 -478 -6195 -472
rect -6129 -438 -6037 -432
rect -6129 -472 -6117 -438
rect -6049 -472 -6037 -438
rect -6129 -478 -6037 -472
rect -5971 -438 -5879 -432
rect -5971 -472 -5959 -438
rect -5891 -472 -5879 -438
rect -5971 -478 -5879 -472
rect -5813 -438 -5721 -432
rect -5813 -472 -5801 -438
rect -5733 -472 -5721 -438
rect -5813 -478 -5721 -472
rect -5655 -438 -5563 -432
rect -5655 -472 -5643 -438
rect -5575 -472 -5563 -438
rect -5655 -478 -5563 -472
rect -5497 -438 -5405 -432
rect -5497 -472 -5485 -438
rect -5417 -472 -5405 -438
rect -5497 -478 -5405 -472
rect -5339 -438 -5247 -432
rect -5339 -472 -5327 -438
rect -5259 -472 -5247 -438
rect -5339 -478 -5247 -472
rect -5181 -438 -5089 -432
rect -5181 -472 -5169 -438
rect -5101 -472 -5089 -438
rect -5181 -478 -5089 -472
rect -5023 -438 -4931 -432
rect -5023 -472 -5011 -438
rect -4943 -472 -4931 -438
rect -5023 -478 -4931 -472
rect -4865 -438 -4773 -432
rect -4865 -472 -4853 -438
rect -4785 -472 -4773 -438
rect -4865 -478 -4773 -472
rect -4707 -438 -4615 -432
rect -4707 -472 -4695 -438
rect -4627 -472 -4615 -438
rect -4707 -478 -4615 -472
rect -4549 -438 -4457 -432
rect -4549 -472 -4537 -438
rect -4469 -472 -4457 -438
rect -4549 -478 -4457 -472
rect -4391 -438 -4299 -432
rect -4391 -472 -4379 -438
rect -4311 -472 -4299 -438
rect -4391 -478 -4299 -472
rect -4233 -438 -4141 -432
rect -4233 -472 -4221 -438
rect -4153 -472 -4141 -438
rect -4233 -478 -4141 -472
rect -4075 -438 -3983 -432
rect -4075 -472 -4063 -438
rect -3995 -472 -3983 -438
rect -4075 -478 -3983 -472
rect -3917 -438 -3825 -432
rect -3917 -472 -3905 -438
rect -3837 -472 -3825 -438
rect -3917 -478 -3825 -472
rect -3759 -438 -3667 -432
rect -3759 -472 -3747 -438
rect -3679 -472 -3667 -438
rect -3759 -478 -3667 -472
rect -3601 -438 -3509 -432
rect -3601 -472 -3589 -438
rect -3521 -472 -3509 -438
rect -3601 -478 -3509 -472
rect -3443 -438 -3351 -432
rect -3443 -472 -3431 -438
rect -3363 -472 -3351 -438
rect -3443 -478 -3351 -472
rect -3285 -438 -3193 -432
rect -3285 -472 -3273 -438
rect -3205 -472 -3193 -438
rect -3285 -478 -3193 -472
rect -3127 -438 -3035 -432
rect -3127 -472 -3115 -438
rect -3047 -472 -3035 -438
rect -3127 -478 -3035 -472
rect -2969 -438 -2877 -432
rect -2969 -472 -2957 -438
rect -2889 -472 -2877 -438
rect -2969 -478 -2877 -472
rect -2811 -438 -2719 -432
rect -2811 -472 -2799 -438
rect -2731 -472 -2719 -438
rect -2811 -478 -2719 -472
rect -2653 -438 -2561 -432
rect -2653 -472 -2641 -438
rect -2573 -472 -2561 -438
rect -2653 -478 -2561 -472
rect -2495 -438 -2403 -432
rect -2495 -472 -2483 -438
rect -2415 -472 -2403 -438
rect -2495 -478 -2403 -472
rect -2337 -438 -2245 -432
rect -2337 -472 -2325 -438
rect -2257 -472 -2245 -438
rect -2337 -478 -2245 -472
rect -2179 -438 -2087 -432
rect -2179 -472 -2167 -438
rect -2099 -472 -2087 -438
rect -2179 -478 -2087 -472
rect -2021 -438 -1929 -432
rect -2021 -472 -2009 -438
rect -1941 -472 -1929 -438
rect -2021 -478 -1929 -472
rect -1863 -438 -1771 -432
rect -1863 -472 -1851 -438
rect -1783 -472 -1771 -438
rect -1863 -478 -1771 -472
rect -1705 -438 -1613 -432
rect -1705 -472 -1693 -438
rect -1625 -472 -1613 -438
rect -1705 -478 -1613 -472
rect -1547 -438 -1455 -432
rect -1547 -472 -1535 -438
rect -1467 -472 -1455 -438
rect -1547 -478 -1455 -472
rect -1389 -438 -1297 -432
rect -1389 -472 -1377 -438
rect -1309 -472 -1297 -438
rect -1389 -478 -1297 -472
rect -1231 -438 -1139 -432
rect -1231 -472 -1219 -438
rect -1151 -472 -1139 -438
rect -1231 -478 -1139 -472
rect -1073 -438 -981 -432
rect -1073 -472 -1061 -438
rect -993 -472 -981 -438
rect -1073 -478 -981 -472
rect -915 -438 -823 -432
rect -915 -472 -903 -438
rect -835 -472 -823 -438
rect -915 -478 -823 -472
rect -757 -438 -665 -432
rect -757 -472 -745 -438
rect -677 -472 -665 -438
rect -757 -478 -665 -472
rect -599 -438 -507 -432
rect -599 -472 -587 -438
rect -519 -472 -507 -438
rect -599 -478 -507 -472
rect -441 -438 -349 -432
rect -441 -472 -429 -438
rect -361 -472 -349 -438
rect -441 -478 -349 -472
rect -283 -438 -191 -432
rect -283 -472 -271 -438
rect -203 -472 -191 -438
rect -283 -478 -191 -472
rect -125 -438 -33 -432
rect -125 -472 -113 -438
rect -45 -472 -33 -438
rect -125 -478 -33 -472
rect 33 -438 125 -432
rect 33 -472 45 -438
rect 113 -472 125 -438
rect 33 -478 125 -472
rect 191 -438 283 -432
rect 191 -472 203 -438
rect 271 -472 283 -438
rect 191 -478 283 -472
rect 349 -438 441 -432
rect 349 -472 361 -438
rect 429 -472 441 -438
rect 349 -478 441 -472
rect 507 -438 599 -432
rect 507 -472 519 -438
rect 587 -472 599 -438
rect 507 -478 599 -472
rect 665 -438 757 -432
rect 665 -472 677 -438
rect 745 -472 757 -438
rect 665 -478 757 -472
rect 823 -438 915 -432
rect 823 -472 835 -438
rect 903 -472 915 -438
rect 823 -478 915 -472
rect 981 -438 1073 -432
rect 981 -472 993 -438
rect 1061 -472 1073 -438
rect 981 -478 1073 -472
rect 1139 -438 1231 -432
rect 1139 -472 1151 -438
rect 1219 -472 1231 -438
rect 1139 -478 1231 -472
rect 1297 -438 1389 -432
rect 1297 -472 1309 -438
rect 1377 -472 1389 -438
rect 1297 -478 1389 -472
rect 1455 -438 1547 -432
rect 1455 -472 1467 -438
rect 1535 -472 1547 -438
rect 1455 -478 1547 -472
rect 1613 -438 1705 -432
rect 1613 -472 1625 -438
rect 1693 -472 1705 -438
rect 1613 -478 1705 -472
rect 1771 -438 1863 -432
rect 1771 -472 1783 -438
rect 1851 -472 1863 -438
rect 1771 -478 1863 -472
rect 1929 -438 2021 -432
rect 1929 -472 1941 -438
rect 2009 -472 2021 -438
rect 1929 -478 2021 -472
rect 2087 -438 2179 -432
rect 2087 -472 2099 -438
rect 2167 -472 2179 -438
rect 2087 -478 2179 -472
rect 2245 -438 2337 -432
rect 2245 -472 2257 -438
rect 2325 -472 2337 -438
rect 2245 -478 2337 -472
rect 2403 -438 2495 -432
rect 2403 -472 2415 -438
rect 2483 -472 2495 -438
rect 2403 -478 2495 -472
rect 2561 -438 2653 -432
rect 2561 -472 2573 -438
rect 2641 -472 2653 -438
rect 2561 -478 2653 -472
rect 2719 -438 2811 -432
rect 2719 -472 2731 -438
rect 2799 -472 2811 -438
rect 2719 -478 2811 -472
rect 2877 -438 2969 -432
rect 2877 -472 2889 -438
rect 2957 -472 2969 -438
rect 2877 -478 2969 -472
rect 3035 -438 3127 -432
rect 3035 -472 3047 -438
rect 3115 -472 3127 -438
rect 3035 -478 3127 -472
rect 3193 -438 3285 -432
rect 3193 -472 3205 -438
rect 3273 -472 3285 -438
rect 3193 -478 3285 -472
rect 3351 -438 3443 -432
rect 3351 -472 3363 -438
rect 3431 -472 3443 -438
rect 3351 -478 3443 -472
rect 3509 -438 3601 -432
rect 3509 -472 3521 -438
rect 3589 -472 3601 -438
rect 3509 -478 3601 -472
rect 3667 -438 3759 -432
rect 3667 -472 3679 -438
rect 3747 -472 3759 -438
rect 3667 -478 3759 -472
rect 3825 -438 3917 -432
rect 3825 -472 3837 -438
rect 3905 -472 3917 -438
rect 3825 -478 3917 -472
rect 3983 -438 4075 -432
rect 3983 -472 3995 -438
rect 4063 -472 4075 -438
rect 3983 -478 4075 -472
rect 4141 -438 4233 -432
rect 4141 -472 4153 -438
rect 4221 -472 4233 -438
rect 4141 -478 4233 -472
rect 4299 -438 4391 -432
rect 4299 -472 4311 -438
rect 4379 -472 4391 -438
rect 4299 -478 4391 -472
rect 4457 -438 4549 -432
rect 4457 -472 4469 -438
rect 4537 -472 4549 -438
rect 4457 -478 4549 -472
rect 4615 -438 4707 -432
rect 4615 -472 4627 -438
rect 4695 -472 4707 -438
rect 4615 -478 4707 -472
rect 4773 -438 4865 -432
rect 4773 -472 4785 -438
rect 4853 -472 4865 -438
rect 4773 -478 4865 -472
rect 4931 -438 5023 -432
rect 4931 -472 4943 -438
rect 5011 -472 5023 -438
rect 4931 -478 5023 -472
rect 5089 -438 5181 -432
rect 5089 -472 5101 -438
rect 5169 -472 5181 -438
rect 5089 -478 5181 -472
rect 5247 -438 5339 -432
rect 5247 -472 5259 -438
rect 5327 -472 5339 -438
rect 5247 -478 5339 -472
rect 5405 -438 5497 -432
rect 5405 -472 5417 -438
rect 5485 -472 5497 -438
rect 5405 -478 5497 -472
rect 5563 -438 5655 -432
rect 5563 -472 5575 -438
rect 5643 -472 5655 -438
rect 5563 -478 5655 -472
rect 5721 -438 5813 -432
rect 5721 -472 5733 -438
rect 5801 -472 5813 -438
rect 5721 -478 5813 -472
rect 5879 -438 5971 -432
rect 5879 -472 5891 -438
rect 5959 -472 5971 -438
rect 5879 -478 5971 -472
rect 6037 -438 6129 -432
rect 6037 -472 6049 -438
rect 6117 -472 6129 -438
rect 6037 -478 6129 -472
rect 6195 -438 6287 -432
rect 6195 -472 6207 -438
rect 6275 -472 6287 -438
rect 6195 -478 6287 -472
<< properties >>
string FIXED_BBOX -6454 -593 6454 593
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.50 m 1 nf 80 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
