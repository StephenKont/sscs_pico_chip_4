magic
tech sky130A
timestamp 1668290293
<< pwell >>
rect -248 -130 248 130
<< nmos >>
rect -150 -25 150 25
<< ndiff >>
rect -179 19 -150 25
rect -179 -19 -173 19
rect -156 -19 -150 19
rect -179 -25 -150 -19
rect 150 19 179 25
rect 150 -19 156 19
rect 173 -19 179 19
rect 150 -25 179 -19
<< ndiffc >>
rect -173 -19 -156 19
rect 156 -19 173 19
<< psubdiff >>
rect -230 95 -182 112
rect 182 95 230 112
rect -230 64 -213 95
rect 213 64 230 95
rect -230 -95 -213 -64
rect 213 -95 230 -64
rect -230 -112 -182 -95
rect 182 -112 230 -95
<< psubdiffcont >>
rect -182 95 182 112
rect -230 -64 -213 64
rect 213 -64 230 64
rect -182 -112 182 -95
<< poly >>
rect -150 61 150 69
rect -150 44 -142 61
rect 142 44 150 61
rect -150 25 150 44
rect -150 -44 150 -25
rect -150 -61 -142 -44
rect 142 -61 150 -44
rect -150 -69 150 -61
<< polycont >>
rect -142 44 142 61
rect -142 -61 142 -44
<< locali >>
rect -230 95 -182 112
rect 182 95 230 112
rect -230 64 -213 95
rect 213 64 230 95
rect -150 44 -142 61
rect 142 44 150 61
rect -173 19 -156 27
rect -173 -27 -156 -19
rect 156 19 173 27
rect 156 -27 173 -19
rect -150 -61 -142 -44
rect 142 -61 150 -44
rect -230 -95 -213 -64
rect 213 -95 230 -64
rect -230 -112 -182 -95
rect 182 -112 230 -95
<< viali >>
rect -142 44 142 61
rect -173 -19 -156 19
rect 156 -19 173 19
rect -142 -61 142 -44
<< metal1 >>
rect -148 61 148 64
rect -148 44 -142 61
rect 142 44 148 61
rect -148 41 148 44
rect -176 19 -153 25
rect -176 -19 -173 19
rect -156 -19 -153 19
rect -176 -25 -153 -19
rect 153 19 176 25
rect 153 -19 156 19
rect 173 -19 176 19
rect 153 -25 176 -19
rect -148 -44 148 -41
rect -148 -61 -142 -44
rect 142 -61 148 -44
rect -148 -64 148 -61
<< properties >>
string FIXED_BBOX -221 -103 221 103
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
