magic
tech sky130A
timestamp 1665559092
<< pwell >>
rect -164 -799 164 799
<< mvnmos >>
rect -50 570 50 670
rect -50 415 50 515
rect -50 260 50 360
rect -50 105 50 205
rect -50 -50 50 50
rect -50 -205 50 -105
rect -50 -360 50 -260
rect -50 -515 50 -415
rect -50 -670 50 -570
<< mvndiff >>
rect -79 664 -50 670
rect -79 576 -73 664
rect -56 576 -50 664
rect -79 570 -50 576
rect 50 664 79 670
rect 50 576 56 664
rect 73 576 79 664
rect 50 570 79 576
rect -79 509 -50 515
rect -79 421 -73 509
rect -56 421 -50 509
rect -79 415 -50 421
rect 50 509 79 515
rect 50 421 56 509
rect 73 421 79 509
rect 50 415 79 421
rect -79 354 -50 360
rect -79 266 -73 354
rect -56 266 -50 354
rect -79 260 -50 266
rect 50 354 79 360
rect 50 266 56 354
rect 73 266 79 354
rect 50 260 79 266
rect -79 199 -50 205
rect -79 111 -73 199
rect -56 111 -50 199
rect -79 105 -50 111
rect 50 199 79 205
rect 50 111 56 199
rect 73 111 79 199
rect 50 105 79 111
rect -79 44 -50 50
rect -79 -44 -73 44
rect -56 -44 -50 44
rect -79 -50 -50 -44
rect 50 44 79 50
rect 50 -44 56 44
rect 73 -44 79 44
rect 50 -50 79 -44
rect -79 -111 -50 -105
rect -79 -199 -73 -111
rect -56 -199 -50 -111
rect -79 -205 -50 -199
rect 50 -111 79 -105
rect 50 -199 56 -111
rect 73 -199 79 -111
rect 50 -205 79 -199
rect -79 -266 -50 -260
rect -79 -354 -73 -266
rect -56 -354 -50 -266
rect -79 -360 -50 -354
rect 50 -266 79 -260
rect 50 -354 56 -266
rect 73 -354 79 -266
rect 50 -360 79 -354
rect -79 -421 -50 -415
rect -79 -509 -73 -421
rect -56 -509 -50 -421
rect -79 -515 -50 -509
rect 50 -421 79 -415
rect 50 -509 56 -421
rect 73 -509 79 -421
rect 50 -515 79 -509
rect -79 -576 -50 -570
rect -79 -664 -73 -576
rect -56 -664 -50 -576
rect -79 -670 -50 -664
rect 50 -576 79 -570
rect 50 -664 56 -576
rect 73 -664 79 -576
rect 50 -670 79 -664
<< mvndiffc >>
rect -73 576 -56 664
rect 56 576 73 664
rect -73 421 -56 509
rect 56 421 73 509
rect -73 266 -56 354
rect 56 266 73 354
rect -73 111 -56 199
rect 56 111 73 199
rect -73 -44 -56 44
rect 56 -44 73 44
rect -73 -199 -56 -111
rect 56 -199 73 -111
rect -73 -354 -56 -266
rect 56 -354 73 -266
rect -73 -509 -56 -421
rect 56 -509 73 -421
rect -73 -664 -56 -576
rect 56 -664 73 -576
<< mvpsubdiff >>
rect -146 775 146 781
rect -146 758 -92 775
rect 92 758 146 775
rect -146 752 146 758
rect -146 727 -117 752
rect -146 -727 -140 727
rect -123 -727 -117 727
rect 117 727 146 752
rect -146 -752 -117 -727
rect 117 -727 123 727
rect 140 -727 146 727
rect 117 -752 146 -727
rect -146 -758 146 -752
rect -146 -775 -92 -758
rect 92 -775 146 -758
rect -146 -781 146 -775
<< mvpsubdiffcont >>
rect -92 758 92 775
rect -140 -727 -123 727
rect 123 -727 140 727
rect -92 -775 92 -758
<< poly >>
rect -50 706 50 714
rect -50 689 -42 706
rect 42 689 50 706
rect -50 670 50 689
rect -50 551 50 570
rect -50 534 -42 551
rect 42 534 50 551
rect -50 515 50 534
rect -50 396 50 415
rect -50 379 -42 396
rect 42 379 50 396
rect -50 360 50 379
rect -50 241 50 260
rect -50 224 -42 241
rect 42 224 50 241
rect -50 205 50 224
rect -50 86 50 105
rect -50 69 -42 86
rect 42 69 50 86
rect -50 50 50 69
rect -50 -69 50 -50
rect -50 -86 -42 -69
rect 42 -86 50 -69
rect -50 -105 50 -86
rect -50 -224 50 -205
rect -50 -241 -42 -224
rect 42 -241 50 -224
rect -50 -260 50 -241
rect -50 -379 50 -360
rect -50 -396 -42 -379
rect 42 -396 50 -379
rect -50 -415 50 -396
rect -50 -534 50 -515
rect -50 -551 -42 -534
rect 42 -551 50 -534
rect -50 -570 50 -551
rect -50 -689 50 -670
rect -50 -706 -42 -689
rect 42 -706 50 -689
rect -50 -714 50 -706
<< polycont >>
rect -42 689 42 706
rect -42 534 42 551
rect -42 379 42 396
rect -42 224 42 241
rect -42 69 42 86
rect -42 -86 42 -69
rect -42 -241 42 -224
rect -42 -396 42 -379
rect -42 -551 42 -534
rect -42 -706 42 -689
<< locali >>
rect -140 758 -92 775
rect 92 758 140 775
rect -140 727 -123 758
rect 123 727 140 758
rect -50 689 -42 706
rect 42 689 50 706
rect -73 664 -56 672
rect -73 568 -56 576
rect 56 664 73 672
rect 56 568 73 576
rect -50 534 -42 551
rect 42 534 50 551
rect -73 509 -56 517
rect -73 413 -56 421
rect 56 509 73 517
rect 56 413 73 421
rect -50 379 -42 396
rect 42 379 50 396
rect -73 354 -56 362
rect -73 258 -56 266
rect 56 354 73 362
rect 56 258 73 266
rect -50 224 -42 241
rect 42 224 50 241
rect -73 199 -56 207
rect -73 103 -56 111
rect 56 199 73 207
rect 56 103 73 111
rect -50 69 -42 86
rect 42 69 50 86
rect -73 44 -56 52
rect -73 -52 -56 -44
rect 56 44 73 52
rect 56 -52 73 -44
rect -50 -86 -42 -69
rect 42 -86 50 -69
rect -73 -111 -56 -103
rect -73 -207 -56 -199
rect 56 -111 73 -103
rect 56 -207 73 -199
rect -50 -241 -42 -224
rect 42 -241 50 -224
rect -73 -266 -56 -258
rect -73 -362 -56 -354
rect 56 -266 73 -258
rect 56 -362 73 -354
rect -50 -396 -42 -379
rect 42 -396 50 -379
rect -73 -421 -56 -413
rect -73 -517 -56 -509
rect 56 -421 73 -413
rect 56 -517 73 -509
rect -50 -551 -42 -534
rect 42 -551 50 -534
rect -73 -576 -56 -568
rect -73 -672 -56 -664
rect 56 -576 73 -568
rect 56 -672 73 -664
rect -50 -706 -42 -689
rect 42 -706 50 -689
rect -140 -758 -123 -727
rect 123 -758 140 -727
rect -140 -775 -92 -758
rect 92 -775 140 -758
<< viali >>
rect -42 689 42 706
rect -73 576 -56 664
rect 56 576 73 664
rect -42 534 42 551
rect -73 421 -56 509
rect 56 421 73 509
rect -42 379 42 396
rect -73 266 -56 354
rect 56 266 73 354
rect -42 224 42 241
rect -73 111 -56 199
rect 56 111 73 199
rect -42 69 42 86
rect -73 -44 -56 44
rect 56 -44 73 44
rect -42 -86 42 -69
rect -73 -199 -56 -111
rect 56 -199 73 -111
rect -42 -241 42 -224
rect -73 -354 -56 -266
rect 56 -354 73 -266
rect -42 -396 42 -379
rect -73 -509 -56 -421
rect 56 -509 73 -421
rect -42 -551 42 -534
rect -73 -664 -56 -576
rect 56 -664 73 -576
rect -42 -706 42 -689
<< metal1 >>
rect -48 706 48 709
rect -48 689 -42 706
rect 42 689 48 706
rect -48 686 48 689
rect -76 664 -53 670
rect -76 576 -73 664
rect -56 576 -53 664
rect -76 570 -53 576
rect 53 664 76 670
rect 53 576 56 664
rect 73 576 76 664
rect 53 570 76 576
rect -48 551 48 554
rect -48 534 -42 551
rect 42 534 48 551
rect -48 531 48 534
rect -76 509 -53 515
rect -76 421 -73 509
rect -56 421 -53 509
rect -76 415 -53 421
rect 53 509 76 515
rect 53 421 56 509
rect 73 421 76 509
rect 53 415 76 421
rect -48 396 48 399
rect -48 379 -42 396
rect 42 379 48 396
rect -48 376 48 379
rect -76 354 -53 360
rect -76 266 -73 354
rect -56 266 -53 354
rect -76 260 -53 266
rect 53 354 76 360
rect 53 266 56 354
rect 73 266 76 354
rect 53 260 76 266
rect -48 241 48 244
rect -48 224 -42 241
rect 42 224 48 241
rect -48 221 48 224
rect -76 199 -53 205
rect -76 111 -73 199
rect -56 111 -53 199
rect -76 105 -53 111
rect 53 199 76 205
rect 53 111 56 199
rect 73 111 76 199
rect 53 105 76 111
rect -48 86 48 89
rect -48 69 -42 86
rect 42 69 48 86
rect -48 66 48 69
rect -76 44 -53 50
rect -76 -44 -73 44
rect -56 -44 -53 44
rect -76 -50 -53 -44
rect 53 44 76 50
rect 53 -44 56 44
rect 73 -44 76 44
rect 53 -50 76 -44
rect -48 -69 48 -66
rect -48 -86 -42 -69
rect 42 -86 48 -69
rect -48 -89 48 -86
rect -76 -111 -53 -105
rect -76 -199 -73 -111
rect -56 -199 -53 -111
rect -76 -205 -53 -199
rect 53 -111 76 -105
rect 53 -199 56 -111
rect 73 -199 76 -111
rect 53 -205 76 -199
rect -48 -224 48 -221
rect -48 -241 -42 -224
rect 42 -241 48 -224
rect -48 -244 48 -241
rect -76 -266 -53 -260
rect -76 -354 -73 -266
rect -56 -354 -53 -266
rect -76 -360 -53 -354
rect 53 -266 76 -260
rect 53 -354 56 -266
rect 73 -354 76 -266
rect 53 -360 76 -354
rect -48 -379 48 -376
rect -48 -396 -42 -379
rect 42 -396 48 -379
rect -48 -399 48 -396
rect -76 -421 -53 -415
rect -76 -509 -73 -421
rect -56 -509 -53 -421
rect -76 -515 -53 -509
rect 53 -421 76 -415
rect 53 -509 56 -421
rect 73 -509 76 -421
rect 53 -515 76 -509
rect -48 -534 48 -531
rect -48 -551 -42 -534
rect 42 -551 48 -534
rect -48 -554 48 -551
rect -76 -576 -53 -570
rect -76 -664 -73 -576
rect -56 -664 -53 -576
rect -76 -670 -53 -664
rect 53 -576 76 -570
rect 53 -664 56 -576
rect 73 -664 76 -576
rect 53 -670 76 -664
rect -48 -689 48 -686
rect -48 -706 -42 -689
rect 42 -706 48 -689
rect -48 -709 48 -706
<< properties >>
string FIXED_BBOX -131 -766 131 766
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 1 m 9 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
