magic
tech sky130A
magscale 1 2
timestamp 1666636516
<< nwell >>
rect -308 -4297 308 4297
<< mvpmos >>
rect -50 -4000 50 4000
<< mvpdiff >>
rect -108 3988 -50 4000
rect -108 -3988 -96 3988
rect -62 -3988 -50 3988
rect -108 -4000 -50 -3988
rect 50 3988 108 4000
rect 50 -3988 62 3988
rect 96 -3988 108 3988
rect 50 -4000 108 -3988
<< mvpdiffc >>
rect -96 -3988 -62 3988
rect 62 -3988 96 3988
<< mvnsubdiff >>
rect -242 4219 242 4231
rect -242 4185 -134 4219
rect 134 4185 242 4219
rect -242 4173 242 4185
rect -242 4123 -184 4173
rect -242 -4123 -230 4123
rect -196 -4123 -184 4123
rect 184 4123 242 4173
rect -242 -4173 -184 -4123
rect 184 -4123 196 4123
rect 230 -4123 242 4123
rect 184 -4173 242 -4123
rect -242 -4185 242 -4173
rect -242 -4219 -134 -4185
rect 134 -4219 242 -4185
rect -242 -4231 242 -4219
<< mvnsubdiffcont >>
rect -134 4185 134 4219
rect -230 -4123 -196 4123
rect 196 -4123 230 4123
rect -134 -4219 134 -4185
<< poly >>
rect -50 4081 50 4097
rect -50 4047 -34 4081
rect 34 4047 50 4081
rect -50 4000 50 4047
rect -50 -4047 50 -4000
rect -50 -4081 -34 -4047
rect 34 -4081 50 -4047
rect -50 -4097 50 -4081
<< polycont >>
rect -34 4047 34 4081
rect -34 -4081 34 -4047
<< locali >>
rect -230 4185 -134 4219
rect 134 4185 230 4219
rect -230 4123 -196 4185
rect 196 4123 230 4185
rect -50 4047 -34 4081
rect 34 4047 50 4081
rect -96 3988 -62 4004
rect -96 -4004 -62 -3988
rect 62 3988 96 4004
rect 62 -4004 96 -3988
rect -50 -4081 -34 -4047
rect 34 -4081 50 -4047
rect -230 -4185 -196 -4123
rect 196 -4185 230 -4123
rect -230 -4219 -134 -4185
rect 134 -4219 230 -4185
<< viali >>
rect -34 4047 34 4081
rect -96 -3988 -62 3988
rect 62 -3988 96 3988
rect -34 -4081 34 -4047
<< metal1 >>
rect -46 4081 46 4087
rect -46 4047 -34 4081
rect 34 4047 46 4081
rect -46 4041 46 4047
rect -102 3988 -56 4000
rect -102 -3988 -96 3988
rect -62 -3988 -56 3988
rect -102 -4000 -56 -3988
rect 56 3988 102 4000
rect 56 -3988 62 3988
rect 96 -3988 102 3988
rect 56 -4000 102 -3988
rect -46 -4047 46 -4041
rect -46 -4081 -34 -4047
rect 34 -4081 46 -4047
rect -46 -4087 46 -4081
<< properties >>
string FIXED_BBOX -213 -4202 213 4202
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 40 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
