magic
tech sky130A
magscale 1 2
timestamp 1667842615
<< viali >>
rect -1282 2672 -1248 2706
rect -854 2666 -820 2700
rect -334 2672 -300 2706
rect 30 2672 64 2706
rect 454 2666 488 2700
rect 688 2672 722 2706
rect 1116 2666 1150 2700
rect 1654 2672 1688 2706
rect 2100 2666 2134 2700
rect 2996 2672 3030 2706
rect 3912 2670 3946 2704
rect 4068 2670 4102 2704
rect 4216 2670 4250 2704
rect 4946 2670 4980 2704
rect 5306 2670 5340 2704
rect 5680 2670 5714 2704
rect 6016 2670 6050 2704
rect 6290 2670 6324 2704
rect 6548 2670 6582 2704
rect 6724 2670 6758 2704
rect 6996 2670 7030 2704
rect 7712 2670 7746 2704
rect 8002 2670 8036 2704
rect 8272 2670 8306 2704
rect 8428 2670 8462 2704
rect 8700 2670 8734 2704
rect 8932 2670 8966 2704
rect 9204 2670 9238 2704
rect 9474 2670 9508 2704
rect 9746 2670 9780 2704
rect 6470 2258 6506 2292
rect 6568 2258 6604 2292
rect 6674 2258 6710 2292
rect 6792 2258 6828 2292
rect 4584 2176 4618 2210
rect 4036 2040 4070 2140
rect 4584 2092 4618 2126
rect 6826 1960 6862 1994
<< metal1 >>
rect 4010 3530 4180 3598
rect -1670 2984 -1616 3034
rect -1628 2980 -1616 2984
rect -1554 2984 -1516 3034
rect -1454 2984 3512 3034
rect 4070 2984 4120 3530
rect 4678 3022 10104 3030
rect -1454 2980 -1438 2984
rect -1628 2972 -1566 2980
rect -1510 2976 -1438 2980
rect -1092 2934 -1056 2984
rect -860 2960 -798 2984
rect -764 2942 -728 2984
rect -436 2944 -400 2984
rect 1206 2940 1242 2984
rect 1532 2944 1568 2984
rect 4678 2980 10010 3022
rect 9982 2968 10010 2980
rect 10072 2968 10104 3022
rect 9982 2950 10104 2968
rect -1758 2874 9942 2924
rect 10226 2816 10276 2842
rect 3646 2814 10276 2816
rect -1670 2768 10276 2814
rect -1670 2766 9870 2768
rect -1288 2706 -1240 2766
rect -1288 2672 -1282 2706
rect -1248 2672 -1240 2706
rect -1288 2660 -1240 2672
rect -862 2700 -814 2766
rect -862 2666 -854 2700
rect -820 2666 -814 2700
rect -862 2654 -814 2666
rect -342 2706 -294 2766
rect -342 2672 -334 2706
rect -300 2672 -294 2706
rect -342 2660 -294 2672
rect 22 2706 70 2766
rect 22 2672 30 2706
rect 64 2672 70 2706
rect 22 2660 70 2672
rect 440 2700 500 2766
rect 440 2666 454 2700
rect 488 2666 500 2700
rect 440 2658 500 2666
rect 680 2706 728 2766
rect 680 2672 688 2706
rect 722 2672 728 2706
rect 680 2660 728 2672
rect 1104 2700 1164 2766
rect 1104 2666 1116 2700
rect 1150 2666 1164 2700
rect 1104 2654 1164 2666
rect 1646 2706 1694 2766
rect 1646 2672 1654 2706
rect 1688 2672 1694 2706
rect 1646 2658 1694 2672
rect 2092 2700 2140 2766
rect 2092 2666 2100 2700
rect 2134 2666 2140 2700
rect 2092 2654 2140 2666
rect 2988 2706 3036 2766
rect 2988 2672 2996 2706
rect 3030 2672 3036 2706
rect 2988 2660 3036 2672
rect 3902 2704 3954 2766
rect 3902 2670 3912 2704
rect 3946 2670 3954 2704
rect 3902 2658 3954 2670
rect 4060 2704 4112 2766
rect 4060 2670 4068 2704
rect 4102 2670 4112 2704
rect 4060 2658 4112 2670
rect 4206 2704 4258 2766
rect 4206 2670 4216 2704
rect 4250 2670 4258 2704
rect 4206 2658 4258 2670
rect 4938 2704 4988 2766
rect 4938 2670 4946 2704
rect 4980 2670 4988 2704
rect 4938 2658 4988 2670
rect 5298 2704 5348 2766
rect 5298 2670 5306 2704
rect 5340 2670 5348 2704
rect 5298 2658 5348 2670
rect 5672 2704 5722 2766
rect 5672 2670 5680 2704
rect 5714 2670 5722 2704
rect 5672 2658 5722 2670
rect 6006 2704 6056 2766
rect 6006 2670 6016 2704
rect 6050 2670 6056 2704
rect 6006 2658 6056 2670
rect 6282 2704 6332 2766
rect 6282 2670 6290 2704
rect 6324 2670 6332 2704
rect 6282 2658 6332 2670
rect 6540 2704 6590 2766
rect 6540 2670 6548 2704
rect 6582 2670 6590 2704
rect 6540 2658 6590 2670
rect 6716 2704 6766 2766
rect 6716 2670 6724 2704
rect 6758 2670 6766 2704
rect 6716 2658 6766 2670
rect 6984 2704 7042 2766
rect 6984 2670 6996 2704
rect 7030 2670 7042 2704
rect 6984 2658 7042 2670
rect 7704 2704 7754 2766
rect 7704 2670 7712 2704
rect 7746 2670 7754 2704
rect 7704 2658 7754 2670
rect 7996 2704 8046 2766
rect 7996 2670 8002 2704
rect 8036 2670 8046 2704
rect 7996 2658 8046 2670
rect 8264 2704 8314 2766
rect 8264 2670 8272 2704
rect 8306 2670 8314 2704
rect 8264 2658 8314 2670
rect 8420 2704 8470 2766
rect 8420 2670 8428 2704
rect 8462 2670 8470 2704
rect 8420 2658 8470 2670
rect 8692 2704 8742 2766
rect 8692 2670 8700 2704
rect 8734 2670 8742 2704
rect 8692 2658 8742 2670
rect 8924 2704 8974 2766
rect 8924 2670 8932 2704
rect 8966 2670 8974 2704
rect 8924 2658 8974 2670
rect 9196 2704 9246 2766
rect 9196 2670 9204 2704
rect 9238 2670 9246 2704
rect 9196 2658 9246 2670
rect 9466 2704 9516 2766
rect 9466 2670 9474 2704
rect 9508 2670 9516 2704
rect 9466 2658 9516 2670
rect 9736 2704 9786 2766
rect 10226 2744 10276 2768
rect 9736 2670 9746 2704
rect 9780 2670 9786 2704
rect 9736 2658 9786 2670
rect 3806 2358 3932 2368
rect 3656 2310 3766 2324
rect 3656 2256 3666 2310
rect 3738 2256 3766 2310
rect 3806 2304 3850 2358
rect 3922 2304 3932 2358
rect 4354 2352 4996 2356
rect 3814 2300 3932 2304
rect 4006 2312 4996 2352
rect 4006 2306 4406 2312
rect 3814 2298 3842 2300
rect 3656 2242 3766 2256
rect 4006 2248 4052 2306
rect 3656 2236 3694 2242
rect 3684 2188 3694 2236
rect 3766 2188 3772 2236
rect 3902 2202 4052 2248
rect 4128 2264 4326 2272
rect 4128 2210 4140 2264
rect 4212 2262 4326 2264
rect 4212 2210 4248 2262
rect 4128 2208 4248 2210
rect 4320 2208 4326 2262
rect 4128 2200 4326 2208
rect 4468 2210 4630 2220
rect 3684 2182 3772 2188
rect 4468 2176 4584 2210
rect 4618 2176 4630 2210
rect 4468 2166 4630 2176
rect 4024 2140 4082 2160
rect 4024 2040 4036 2140
rect 4070 2040 4082 2140
rect 4024 1942 4082 2040
rect 4466 2126 4630 2134
rect 4466 2092 4584 2126
rect 4618 2092 4630 2126
rect 4466 2082 4630 2092
rect 4934 2090 4996 2312
rect 6450 2292 6520 2314
rect 6450 2258 6470 2292
rect 6506 2258 6520 2292
rect 6450 2094 6520 2258
rect 6552 2292 6622 2312
rect 6552 2258 6568 2292
rect 6604 2258 6622 2292
rect 6552 2092 6622 2258
rect 6658 2292 6728 2312
rect 6658 2258 6674 2292
rect 6710 2258 6728 2292
rect 6658 2092 6728 2258
rect 6774 2292 6844 2312
rect 6774 2258 6792 2292
rect 6828 2258 6844 2292
rect 6774 2162 6844 2258
rect 6774 2092 6876 2162
rect 4466 1944 4512 2082
rect 6814 1994 6876 2092
rect 6814 1960 6826 1994
rect 6862 1960 6876 1994
rect 6814 1944 6876 1960
rect 4466 1942 6876 1944
rect 4024 1896 6876 1942
<< via1 >>
rect -1616 2980 -1554 3034
rect -1516 2980 -1454 3034
rect 10010 2968 10072 3022
rect 3666 2256 3738 2310
rect 3850 2304 3922 2358
rect 3694 2188 3766 2242
rect 4140 2210 4212 2264
rect 4248 2208 4320 2262
<< metal2 >>
rect -1890 3034 -1438 3036
rect -1890 2980 -1616 3034
rect -1554 2980 -1516 3034
rect -1454 2980 -1438 3034
rect -1890 2968 -1438 2980
rect -1890 2324 -1810 2968
rect -1518 2956 -1438 2968
rect 9982 3022 10104 3030
rect 9982 2968 10010 3022
rect 10072 2968 10104 3022
rect 9982 2950 10104 2968
rect 10036 2494 10104 2950
rect 4240 2426 10104 2494
rect 3806 2358 3932 2370
rect -1890 2316 3772 2324
rect -1888 2310 3772 2316
rect -1888 2256 3666 2310
rect 3738 2256 3772 2310
rect 3806 2304 3850 2358
rect 3922 2356 3932 2358
rect 4240 2356 4308 2426
rect 3922 2320 4326 2356
rect 3922 2304 3932 2320
rect 3806 2300 3932 2304
rect -1888 2242 3772 2256
rect -1888 2236 3694 2242
rect 3684 2188 3694 2236
rect 3766 2188 3772 2242
rect 4128 2264 4326 2320
rect 4128 2210 4140 2264
rect 4212 2262 4326 2264
rect 4212 2210 4248 2262
rect 4128 2208 4248 2210
rect 4320 2208 4326 2262
rect 4128 2200 4326 2208
rect 3684 2182 3772 2188
use sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ  sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ_0
timestamp 1666571082
transform 1 0 3840 0 1 2172
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ  sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ_1
timestamp 1666571082
transform 1 0 4388 0 1 2168
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_5FQFS2  sky130_fd_pr__pfet_g5v0d10v5_5FQFS2_0
timestamp 1665420977
transform 0 1 7295 -1 0 2900
box -308 -2857 308 2857
use sky130_fd_pr__pfet_g5v0d10v5_5FQFS2  sky130_fd_pr__pfet_g5v0d10v5_5FQFS2_1
timestamp 1665420977
transform 0 1 895 -1 0 2902
box -308 -2857 308 2857
use sky130_fd_pr__pfet_g5v0d10v5_AJQB7U  sky130_fd_pr__pfet_g5v0d10v5_AJQB7U_0
timestamp 1666571082
transform 0 1 4095 1 0 2900
box -308 -397 308 397
use sky130_fd_pr__res_high_po_0p35_MTJUHY  sky130_fd_pr__res_high_po_0p35_MTJUHY_0
timestamp 1665495179
transform 0 1 5889 -1 0 2127
box -201 -1133 201 1133
<< labels >>
rlabel metal1 10226 2744 10276 2842 1 Vdd
port 2 n
rlabel metal1 4010 3530 4180 3598 1 out_current
port 1 n
<< end >>
