magic
tech sky130A
magscale 1 2
timestamp 1665942722
<< error_p >>
rect -287 225 -225 231
rect -159 225 -97 231
rect -31 225 31 231
rect 97 225 159 231
rect 225 225 287 231
rect -287 191 -275 225
rect -159 191 -147 225
rect -31 191 -19 225
rect 97 191 109 225
rect 225 191 237 225
rect -287 185 -225 191
rect -159 185 -97 191
rect -31 185 31 191
rect 97 185 159 191
rect 225 185 287 191
rect -287 -191 -225 -185
rect -159 -191 -97 -185
rect -31 -191 31 -185
rect 97 -191 159 -185
rect 225 -191 287 -185
rect -287 -225 -275 -191
rect -159 -225 -147 -191
rect -31 -225 -19 -191
rect 97 -225 109 -191
rect 225 -225 237 -191
rect -287 -231 -225 -225
rect -159 -231 -97 -225
rect -31 -231 31 -225
rect 97 -231 159 -225
rect 225 -231 287 -225
<< nwell >>
rect -487 -363 487 363
<< pmoslvt >>
rect -291 -144 -221 144
rect -163 -144 -93 144
rect -35 -144 35 144
rect 93 -144 163 144
rect 221 -144 291 144
<< pdiff >>
rect -349 132 -291 144
rect -349 -132 -337 132
rect -303 -132 -291 132
rect -349 -144 -291 -132
rect -221 132 -163 144
rect -221 -132 -209 132
rect -175 -132 -163 132
rect -221 -144 -163 -132
rect -93 132 -35 144
rect -93 -132 -81 132
rect -47 -132 -35 132
rect -93 -144 -35 -132
rect 35 132 93 144
rect 35 -132 47 132
rect 81 -132 93 132
rect 35 -144 93 -132
rect 163 132 221 144
rect 163 -132 175 132
rect 209 -132 221 132
rect 163 -144 221 -132
rect 291 132 349 144
rect 291 -132 303 132
rect 337 -132 349 132
rect 291 -144 349 -132
<< pdiffc >>
rect -337 -132 -303 132
rect -209 -132 -175 132
rect -81 -132 -47 132
rect 47 -132 81 132
rect 175 -132 209 132
rect 303 -132 337 132
<< nsubdiff >>
rect -451 293 -355 327
rect 355 293 451 327
rect -451 231 -417 293
rect 417 231 451 293
rect -451 -293 -417 -231
rect 417 -293 451 -231
rect -451 -327 -355 -293
rect 355 -327 451 -293
<< nsubdiffcont >>
rect -355 293 355 327
rect -451 -231 -417 231
rect 417 -231 451 231
rect -355 -327 355 -293
<< poly >>
rect -291 225 -221 241
rect -291 191 -275 225
rect -237 191 -221 225
rect -291 144 -221 191
rect -163 225 -93 241
rect -163 191 -147 225
rect -109 191 -93 225
rect -163 144 -93 191
rect -35 225 35 241
rect -35 191 -19 225
rect 19 191 35 225
rect -35 144 35 191
rect 93 225 163 241
rect 93 191 109 225
rect 147 191 163 225
rect 93 144 163 191
rect 221 225 291 241
rect 221 191 237 225
rect 275 191 291 225
rect 221 144 291 191
rect -291 -191 -221 -144
rect -291 -225 -275 -191
rect -237 -225 -221 -191
rect -291 -241 -221 -225
rect -163 -191 -93 -144
rect -163 -225 -147 -191
rect -109 -225 -93 -191
rect -163 -241 -93 -225
rect -35 -191 35 -144
rect -35 -225 -19 -191
rect 19 -225 35 -191
rect -35 -241 35 -225
rect 93 -191 163 -144
rect 93 -225 109 -191
rect 147 -225 163 -191
rect 93 -241 163 -225
rect 221 -191 291 -144
rect 221 -225 237 -191
rect 275 -225 291 -191
rect 221 -241 291 -225
<< polycont >>
rect -275 191 -237 225
rect -147 191 -109 225
rect -19 191 19 225
rect 109 191 147 225
rect 237 191 275 225
rect -275 -225 -237 -191
rect -147 -225 -109 -191
rect -19 -225 19 -191
rect 109 -225 147 -191
rect 237 -225 275 -191
<< locali >>
rect -451 293 -355 327
rect 355 293 451 327
rect -451 231 -417 293
rect 417 231 451 293
rect -291 191 -275 225
rect -237 191 -221 225
rect -163 191 -147 225
rect -109 191 -93 225
rect -35 191 -19 225
rect 19 191 35 225
rect 93 191 109 225
rect 147 191 163 225
rect 221 191 237 225
rect 275 191 291 225
rect -337 132 -303 148
rect -337 -148 -303 -132
rect -209 132 -175 148
rect -209 -148 -175 -132
rect -81 132 -47 148
rect -81 -148 -47 -132
rect 47 132 81 148
rect 47 -148 81 -132
rect 175 132 209 148
rect 175 -148 209 -132
rect 303 132 337 148
rect 303 -148 337 -132
rect -291 -225 -275 -191
rect -237 -225 -221 -191
rect -163 -225 -147 -191
rect -109 -225 -93 -191
rect -35 -225 -19 -191
rect 19 -225 35 -191
rect 93 -225 109 -191
rect 147 -225 163 -191
rect 221 -225 237 -191
rect 275 -225 291 -191
rect -451 -293 -417 -231
rect 417 -293 451 -231
rect -451 -327 -355 -293
rect 355 -327 451 -293
<< viali >>
rect -275 191 -237 225
rect -147 191 -109 225
rect -19 191 19 225
rect 109 191 147 225
rect 237 191 275 225
rect -337 -132 -303 132
rect -209 -132 -175 132
rect -81 -132 -47 132
rect 47 -132 81 132
rect 175 -132 209 132
rect 303 -132 337 132
rect -275 -225 -237 -191
rect -147 -225 -109 -191
rect -19 -225 19 -191
rect 109 -225 147 -191
rect 237 -225 275 -191
<< metal1 >>
rect -287 225 -225 231
rect -287 191 -275 225
rect -237 191 -225 225
rect -287 185 -225 191
rect -159 225 -97 231
rect -159 191 -147 225
rect -109 191 -97 225
rect -159 185 -97 191
rect -31 225 31 231
rect -31 191 -19 225
rect 19 191 31 225
rect -31 185 31 191
rect 97 225 159 231
rect 97 191 109 225
rect 147 191 159 225
rect 97 185 159 191
rect 225 225 287 231
rect 225 191 237 225
rect 275 191 287 225
rect 225 185 287 191
rect -343 132 -297 144
rect -343 -132 -337 132
rect -303 -132 -297 132
rect -343 -144 -297 -132
rect -215 132 -169 144
rect -215 -132 -209 132
rect -175 -132 -169 132
rect -215 -144 -169 -132
rect -87 132 -41 144
rect -87 -132 -81 132
rect -47 -132 -41 132
rect -87 -144 -41 -132
rect 41 132 87 144
rect 41 -132 47 132
rect 81 -132 87 132
rect 41 -144 87 -132
rect 169 132 215 144
rect 169 -132 175 132
rect 209 -132 215 132
rect 169 -144 215 -132
rect 297 132 343 144
rect 297 -132 303 132
rect 337 -132 343 132
rect 297 -144 343 -132
rect -287 -191 -225 -185
rect -287 -225 -275 -191
rect -237 -225 -225 -191
rect -287 -231 -225 -225
rect -159 -191 -97 -185
rect -159 -225 -147 -191
rect -109 -225 -97 -191
rect -159 -231 -97 -225
rect -31 -191 31 -185
rect -31 -225 -19 -191
rect 19 -225 31 -191
rect -31 -231 31 -225
rect 97 -191 159 -185
rect 97 -225 109 -191
rect 147 -225 159 -191
rect 97 -231 159 -225
rect 225 -191 287 -185
rect 225 -225 237 -191
rect 275 -225 287 -191
rect 225 -231 287 -225
<< properties >>
string FIXED_BBOX -434 -310 434 310
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.44 l 0.35 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
