magic
tech sky130A
magscale 1 2
timestamp 1667842615
<< nwell >>
rect 11468 255 11546 627
<< pwell >>
rect 11429 -28 11589 2
rect 11426 -77 11589 -28
<< locali >>
rect 3480 1194 3636 1244
rect 6264 1198 6420 1244
rect 8856 1194 9012 1244
rect 3480 600 3636 650
rect 6264 602 6420 648
rect 8856 600 9012 650
rect 24 526 180 582
rect 11399 572 11732 606
rect 11602 524 11758 572
rect 649 123 703 359
rect 24 -62 180 -14
rect 11602 -60 11758 -14
rect 2520 -134 2676 -76
rect 5208 -132 5364 -86
rect 7992 -132 8148 -80
rect 10776 -136 10932 -72
rect 11303 -94 11758 -60
rect 2520 -732 2676 -674
rect 5208 -728 5364 -682
rect 7992 -732 8148 -680
rect 2040 -800 2196 -738
rect 3864 -804 4020 -740
rect 10776 -742 10932 -678
rect 4728 -800 4884 -746
rect 6552 -808 6708 -754
rect 7416 -810 7572 -754
rect 9240 -802 9396 -746
rect 10104 -802 10260 -744
rect 11928 -802 12084 -750
rect 2040 -1402 2196 -1340
rect 3864 -1396 4020 -1332
rect 4728 -1398 4884 -1344
rect 6552 -1398 6708 -1344
rect 7416 -1400 7572 -1344
rect 9240 -1400 9396 -1344
rect 10104 -1398 10260 -1340
rect 11928 -1400 12084 -1348
rect 2904 -1468 3060 -1422
rect 5592 -1468 5748 -1422
rect 8184 -1468 8340 -1422
rect 10872 -1468 11028 -1422
rect 2904 -2062 3060 -2016
rect 5592 -2062 5748 -2016
rect 8184 -2064 8340 -2018
rect 10872 -2060 11028 -2014
rect 2346 -4333 2802 -4299
rect 2919 -4333 3376 -4299
rect 1227 -6743 1367 -6709
rect 2798 -6725 2924 -6691
rect 2346 -18333 2802 -18299
rect 2919 -18333 3376 -18299
rect 1227 -20743 1367 -20709
rect 2798 -20725 2924 -20691
rect 2346 -32333 2802 -32299
rect 2919 -32333 3376 -32299
rect 1227 -34743 1367 -34709
rect 2798 -34725 2924 -34691
rect 2346 -46333 2802 -46299
rect 2919 -46333 3376 -46299
rect 1227 -48743 1367 -48709
rect 2798 -48725 2924 -48691
<< viali >>
rect 219 159 294 233
rect 401 167 467 233
rect 511 159 581 233
rect 3589 313 3623 347
rect 6277 313 6311 347
rect 8965 313 8999 347
rect 892 165 926 267
rect 1068 185 1133 251
rect 3298 177 3392 279
rect 3580 165 3614 267
rect 3756 185 3821 251
rect 5986 177 6080 279
rect 6268 165 6302 267
rect 6444 185 6509 251
rect 8674 177 8768 279
rect 8956 165 8990 267
rect 9132 185 9197 251
rect 11362 177 11456 279
rect 19112 -423 19380 -389
rect 19016 -931 19050 -485
rect 19442 -931 19476 -485
rect 19112 -1027 19380 -993
rect 19124 -1281 19392 -1247
rect 19028 -1771 19062 -1343
rect 19454 -1771 19488 -1343
rect 19124 -1867 19392 -1833
rect 11516 -2470 12778 -2436
rect 13046 -2470 14308 -2436
rect 11420 -2670 11454 -2532
rect 12840 -2670 12874 -2532
rect 12950 -2670 12984 -2532
rect 14370 -2670 14404 -2532
rect 11516 -2766 12778 -2732
rect 13046 -2766 14308 -2732
rect 630 -3719 1980 -3685
rect 534 -4955 568 -3874
rect 2042 -4955 2076 -3781
rect 2250 -4951 2284 -4395
rect 3438 -4951 3472 -4395
rect 630 -5051 1980 -5017
rect 2346 -5047 3376 -5013
rect 630 -5411 1980 -5377
rect 534 -6647 568 -5473
rect 2042 -6647 2076 -5473
rect 2346 -6211 2621 -6177
rect 3101 -6211 3376 -6177
rect 2250 -6629 2284 -6273
rect 3438 -6629 3472 -6273
rect 630 -6743 1221 -6709
rect 1373 -6743 1980 -6709
rect 2346 -6725 2792 -6691
rect 2930 -6725 3376 -6691
rect 41068 -11777 42114 -11743
rect 630 -17719 1980 -17685
rect 534 -18955 568 -17874
rect 2042 -18955 2076 -17781
rect 2250 -18951 2284 -18395
rect 3438 -18951 3472 -18395
rect 630 -19051 1980 -19017
rect 2346 -19047 3376 -19013
rect 630 -19411 1980 -19377
rect 534 -20647 568 -19473
rect 2042 -20647 2076 -19473
rect 2346 -20211 2621 -20177
rect 3101 -20211 3376 -20177
rect 2250 -20629 2284 -20273
rect 3438 -20629 3472 -20273
rect 630 -20743 1221 -20709
rect 1373 -20743 1980 -20709
rect 2346 -20725 2792 -20691
rect 2930 -20725 3376 -20691
rect 40972 -24589 41006 -11839
rect 42176 -24589 42210 -11839
rect 41068 -24685 42114 -24651
rect 630 -31719 1980 -31685
rect 534 -32955 568 -31874
rect 2042 -32955 2076 -31781
rect 2250 -32951 2284 -32395
rect 3438 -32951 3472 -32395
rect 630 -33051 1980 -33017
rect 2346 -33047 3376 -33013
rect 630 -33411 1980 -33377
rect 534 -34647 568 -33473
rect 2042 -34647 2076 -33473
rect 2346 -34211 2621 -34177
rect 3101 -34211 3376 -34177
rect 2250 -34629 2284 -34273
rect 3438 -34629 3472 -34273
rect 630 -34743 1221 -34709
rect 1373 -34743 1980 -34709
rect 2346 -34725 2792 -34691
rect 2930 -34725 3376 -34691
rect 630 -45719 1980 -45685
rect 534 -46955 568 -45874
rect 2042 -46955 2076 -45781
rect 2250 -46951 2284 -46395
rect 3438 -46951 3472 -46395
rect 630 -47051 1980 -47017
rect 2346 -47047 3376 -47013
rect 630 -47411 1980 -47377
rect 534 -48647 568 -47473
rect 2042 -48647 2076 -47473
rect 2346 -48211 2621 -48177
rect 3101 -48211 3376 -48177
rect 2250 -48629 2284 -48273
rect 3438 -48629 3472 -48273
rect 630 -48743 1221 -48709
rect 1373 -48743 1980 -48709
rect 2346 -48725 2792 -48691
rect 2930 -48725 3376 -48691
<< metal1 >>
rect -607 1206 9190 1304
rect -607 -28 -268 1206
rect 12540 831 12928 983
rect 12540 739 12686 831
rect 12778 739 12928 831
rect -196 638 -98 644
rect -98 540 11674 638
rect 12540 586 12928 739
rect 19038 720 19500 784
rect -196 534 -98 540
rect 879 346 947 353
rect 501 259 614 267
rect 371 246 473 252
rect 205 239 303 245
rect 205 153 211 239
rect 297 153 303 239
rect 371 160 377 246
rect 467 160 473 246
rect 371 154 473 160
rect 501 233 517 259
rect 501 159 511 233
rect 607 165 614 259
rect 581 159 614 165
rect 205 147 303 153
rect 501 147 614 159
rect 879 162 885 346
rect 937 162 947 346
rect 3567 347 3635 353
rect 3567 346 3589 347
rect 3623 346 3635 347
rect 3286 279 3404 291
rect 1056 257 1145 263
rect 1056 179 1062 257
rect 1137 179 1145 257
rect 1056 173 1145 179
rect 3286 177 3298 279
rect 3392 177 3404 279
rect 3286 165 3404 177
rect 879 156 947 162
rect 3567 162 3573 346
rect 3625 162 3635 346
rect 6255 347 6323 353
rect 6255 346 6277 347
rect 6311 346 6323 347
rect 5975 279 6092 291
rect 3744 257 3833 263
rect 3744 179 3750 257
rect 3825 179 3833 257
rect 3744 173 3833 179
rect 5975 177 5986 279
rect 6080 177 6092 279
rect 5975 165 6092 177
rect 3567 156 3635 162
rect 6255 162 6261 346
rect 6313 162 6323 346
rect 8943 347 9011 353
rect 8943 346 8965 347
rect 8999 346 9011 347
rect 8663 279 8780 291
rect 6432 257 6521 263
rect 6432 179 6438 257
rect 6513 179 6521 257
rect 6432 173 6521 179
rect 8663 177 8674 279
rect 8768 177 8780 279
rect 8663 165 8780 177
rect 6255 156 6323 162
rect 8943 162 8949 346
rect 9001 162 9011 346
rect 11351 279 11468 291
rect 9120 257 9209 263
rect 9120 179 9126 257
rect 9201 179 9209 257
rect 9120 173 9209 179
rect 11351 177 11362 279
rect 11456 177 11468 279
rect 11351 165 11468 177
rect 8943 156 9011 162
rect -6127 -213 -5411 -70
rect -607 -126 11674 -28
rect -607 -213 -268 -126
rect -6127 -552 -5966 -213
rect -5627 -552 -267 -213
rect -6127 -683 -5411 -552
rect -607 -1360 -268 -552
rect -196 -694 -98 -688
rect -98 -792 11674 -694
rect -196 -798 -98 -792
rect 2599 -893 2883 -879
rect 2599 -1012 2615 -893
rect 2865 -1012 2883 -893
rect 2599 -1025 2883 -1012
rect 5287 -893 5571 -879
rect 5287 -1002 5303 -893
rect 5553 -1002 5571 -893
rect 5287 -1025 5571 -1002
rect 7975 -903 8259 -879
rect 7975 -1007 8001 -903
rect 8222 -1007 8259 -903
rect 7975 -1025 8259 -1007
rect 10663 -903 10947 -879
rect 10663 -1006 10686 -903
rect 10902 -1006 10947 -903
rect 10663 -1025 10947 -1006
rect 3292 -1058 3576 -1053
rect 3292 -1189 3298 -1058
rect 3565 -1189 3576 -1058
rect 8668 -1072 8952 -1053
rect 3292 -1199 3576 -1189
rect 5980 -1189 5986 -1078
rect 6253 -1189 6264 -1078
rect 8668 -1159 8692 -1072
rect 8926 -1159 8952 -1072
rect 8668 -1172 8952 -1159
rect 11356 -1078 11640 -1053
rect 11356 -1166 11378 -1078
rect 11608 -1166 11640 -1078
rect 11356 -1182 11640 -1166
rect 5980 -1199 6264 -1189
rect 12686 -1266 12778 586
rect 19038 400 19140 720
rect 19460 661 19500 720
rect 19460 489 41568 661
rect 19460 400 19500 489
rect 19038 337 19500 400
rect 19160 52 19437 67
rect 19160 -206 19171 52
rect 19429 -206 19437 52
rect 19160 -216 19437 -206
rect 19203 -376 19381 -216
rect 19003 -389 19488 -376
rect 19003 -423 19112 -389
rect 19380 -423 19488 -389
rect 19003 -435 19488 -423
rect 19003 -485 19062 -435
rect 19003 -931 19016 -485
rect 19050 -608 19062 -485
rect 19429 -485 19488 -435
rect 19050 -808 19190 -608
rect 19296 -615 19365 -608
rect 19296 -802 19302 -615
rect 19354 -802 19365 -615
rect 19296 -808 19365 -802
rect 19050 -931 19062 -808
rect 19003 -980 19062 -931
rect 19196 -862 19296 -849
rect 19196 -933 19206 -862
rect 19286 -933 19296 -862
rect 19196 -943 19296 -933
rect 19429 -931 19442 -485
rect 19476 -931 19488 -485
rect 19429 -980 19488 -931
rect 19003 -993 19488 -980
rect 19003 -1027 19112 -993
rect 19380 -1027 19488 -993
rect 19003 -1039 19488 -1027
rect 12866 -1149 13076 -1132
rect 12866 -1219 12873 -1149
rect 12943 -1219 13076 -1149
rect 12866 -1222 13076 -1219
rect 19016 -1247 19500 -1235
rect 12686 -1358 13074 -1266
rect 19016 -1281 19124 -1247
rect 19392 -1281 19500 -1247
rect 19016 -1293 19500 -1281
rect 19016 -1343 19074 -1293
rect -607 -1458 12026 -1360
rect 18769 -1483 18951 -1471
rect 19016 -1483 19028 -1343
rect 18769 -1648 18779 -1483
rect 18944 -1648 19028 -1483
rect 18769 -1654 18951 -1648
rect 19016 -1771 19028 -1648
rect 19062 -1457 19074 -1343
rect 19208 -1347 19308 -1336
rect 19208 -1414 19217 -1347
rect 19298 -1414 19308 -1347
rect 19208 -1425 19308 -1414
rect 19442 -1343 19500 -1293
rect 19062 -1657 19201 -1457
rect 19308 -1466 19374 -1457
rect 19308 -1650 19315 -1466
rect 19367 -1650 19374 -1466
rect 19308 -1657 19374 -1650
rect 19062 -1771 19074 -1657
rect 19016 -1821 19074 -1771
rect 19442 -1771 19454 -1343
rect 19488 -1771 19500 -1343
rect 19442 -1821 19500 -1771
rect 19016 -1833 19500 -1821
rect 19016 -1867 19124 -1833
rect 19392 -1867 19500 -1833
rect 19016 -1879 19500 -1867
rect -202 -2124 -196 -2026
rect -98 -2124 11298 -2026
rect 14181 -2133 14187 -2043
rect 14277 -2133 14283 -2043
rect 14187 -2400 14277 -2133
rect 2593 -2710 2599 -2426
rect 2883 -2710 2889 -2426
rect 5281 -2710 5287 -2426
rect 5571 -2710 5577 -2426
rect 7969 -2710 7975 -2426
rect 8259 -2710 8265 -2426
rect 10657 -2710 10663 -2426
rect 10947 -2710 10953 -2426
rect 11384 -2436 14440 -2400
rect 11384 -2470 11516 -2436
rect 12778 -2470 13046 -2436
rect 14308 -2470 14440 -2436
rect 11384 -2490 14440 -2470
rect 11384 -2532 11474 -2490
rect 11384 -2670 11420 -2532
rect 11454 -2670 11474 -2532
rect 11550 -2636 11982 -2490
rect 12820 -2532 13004 -2490
rect 12312 -2572 12744 -2566
rect 12312 -2630 12320 -2572
rect 12736 -2630 12744 -2572
rect 12312 -2636 12744 -2630
rect 2599 -3524 2883 -2710
rect 3286 -3290 3292 -3006
rect 3576 -3290 4056 -3006
rect 368 -3580 3619 -3524
rect 368 -3771 424 -3580
rect 606 -3656 2112 -3649
rect 606 -3685 642 -3656
rect 1967 -3685 2112 -3656
rect 606 -3719 630 -3685
rect 1980 -3719 2112 -3685
rect 606 -3729 642 -3719
rect 1967 -3729 2112 -3719
rect 606 -3735 2112 -3729
rect 368 -3827 822 -3771
rect 2022 -3781 2112 -3735
rect 368 -4898 424 -3827
rect 2022 -3868 2042 -3781
rect 498 -3874 694 -3868
rect 360 -4912 432 -4898
rect 360 -4968 368 -4912
rect 424 -4968 432 -4912
rect 360 -4974 432 -4968
rect 498 -4955 534 -3874
rect 568 -3875 694 -3874
rect 568 -4862 639 -3875
rect 692 -4862 694 -3875
rect 568 -4868 694 -4862
rect 764 -3875 822 -3868
rect 764 -4862 767 -3875
rect 820 -4862 822 -3875
rect 764 -4868 822 -4862
rect 892 -3875 950 -3868
rect 892 -4862 895 -3875
rect 948 -4862 950 -3875
rect 892 -4868 950 -4862
rect 1020 -3875 1078 -3868
rect 1020 -4862 1023 -3875
rect 1076 -4862 1078 -3875
rect 1020 -4868 1078 -4862
rect 1148 -3875 1206 -3868
rect 1148 -4862 1151 -3875
rect 1204 -4862 1206 -3875
rect 1148 -4868 1206 -4862
rect 1276 -3875 1334 -3868
rect 1276 -4862 1279 -3875
rect 1332 -4862 1334 -3875
rect 1276 -4868 1334 -4862
rect 1404 -3875 1462 -3868
rect 1404 -4862 1407 -3875
rect 1460 -4862 1462 -3875
rect 1404 -4868 1462 -4862
rect 1532 -3875 1590 -3868
rect 1532 -4862 1535 -3875
rect 1588 -4862 1590 -3875
rect 1532 -4868 1590 -4862
rect 1660 -3875 1718 -3868
rect 1660 -4862 1663 -3875
rect 1716 -4862 1718 -3875
rect 1660 -4868 1718 -4862
rect 1788 -3875 1846 -3868
rect 1788 -4862 1791 -3875
rect 1844 -4862 1846 -3875
rect 1788 -4868 1846 -4862
rect 1916 -3875 2042 -3868
rect 1916 -4862 1919 -3875
rect 1972 -4862 2042 -3875
rect 1916 -4868 2042 -4862
rect 568 -4955 578 -4868
rect 498 -5008 578 -4955
rect 614 -4909 682 -4903
rect 1904 -4907 1989 -4901
rect 1904 -4909 1911 -4907
rect 614 -4965 620 -4909
rect 676 -4965 946 -4909
rect 1896 -4960 1911 -4909
rect 1983 -4960 1989 -4907
rect 1896 -4965 1989 -4960
rect 2022 -4955 2042 -4868
rect 2076 -4955 2112 -3781
rect 614 -4971 682 -4965
rect 2022 -5008 2112 -4955
rect 498 -5017 2112 -5008
rect 498 -5051 630 -5017
rect 1980 -5051 2112 -5017
rect 498 -5087 2112 -5051
rect 498 -5341 602 -5087
rect 2008 -5341 2112 -5087
rect 498 -5377 2112 -5341
rect 498 -5411 630 -5377
rect 1980 -5411 2112 -5377
rect 498 -5427 2112 -5411
rect 498 -5473 588 -5427
rect 498 -6647 534 -5473
rect 568 -6647 588 -5473
rect 1902 -5461 1987 -5455
rect 1902 -5514 1909 -5461
rect 1981 -5514 1987 -5461
rect 1902 -5519 1987 -5514
rect 2022 -5473 2112 -5427
rect 636 -5567 694 -5560
rect 636 -6554 639 -5567
rect 692 -6554 694 -5567
rect 636 -6560 694 -6554
rect 764 -5567 822 -5560
rect 764 -6554 767 -5567
rect 820 -6554 822 -5567
rect 764 -6560 822 -6554
rect 892 -5567 950 -5560
rect 892 -6554 895 -5567
rect 948 -6554 950 -5567
rect 892 -6560 950 -6554
rect 1020 -5567 1078 -5560
rect 1020 -6554 1023 -5567
rect 1076 -6554 1078 -5567
rect 1020 -6560 1078 -6554
rect 1148 -5567 1206 -5560
rect 1148 -6554 1151 -5567
rect 1204 -6554 1206 -5567
rect 1148 -6560 1206 -6554
rect 1276 -5567 1334 -5560
rect 1276 -6554 1279 -5567
rect 1332 -6554 1334 -5567
rect 1276 -6560 1334 -6554
rect 1404 -5567 1462 -5560
rect 1404 -6554 1407 -5567
rect 1460 -6554 1462 -5567
rect 1404 -6560 1462 -6554
rect 1532 -5567 1590 -5560
rect 1532 -6554 1535 -5567
rect 1588 -6554 1590 -5567
rect 1532 -6560 1590 -6554
rect 1660 -5567 1718 -5560
rect 1660 -6554 1663 -5567
rect 1716 -6554 1718 -5567
rect 1660 -6560 1718 -6554
rect 1788 -5567 1846 -5560
rect 1788 -6554 1791 -5567
rect 1844 -6554 1846 -5567
rect 1788 -6560 1846 -6554
rect 1916 -5567 1974 -5560
rect 1916 -6554 1919 -5567
rect 1972 -6554 1974 -5567
rect 1916 -6560 1974 -6554
rect 498 -6693 588 -6647
rect 498 -6709 1227 -6693
rect 498 -6743 630 -6709
rect 1221 -6743 1227 -6709
rect 498 -6779 1227 -6743
rect 1269 -6822 1339 -6629
rect 2022 -6647 2042 -5473
rect 2076 -6647 2112 -5473
rect 2022 -6693 2112 -6647
rect 1367 -6709 2112 -6693
rect 1367 -6743 1373 -6709
rect 1980 -6743 2112 -6709
rect 1367 -6779 2112 -6743
rect 2214 -4340 2802 -4263
rect 2214 -4395 2304 -4340
rect 2834 -4385 2890 -3580
rect 3563 -3863 3619 -3580
rect 3541 -3888 3646 -3863
rect 3541 -3944 3563 -3888
rect 3619 -3944 3646 -3888
rect 3541 -3961 3646 -3944
rect 2919 -4340 3508 -4263
rect 2214 -4951 2250 -4395
rect 2284 -4951 2304 -4395
rect 2492 -4441 3326 -4385
rect 3432 -4395 3508 -4340
rect 2348 -4867 2354 -4473
rect 2408 -4867 2414 -4473
rect 2348 -4873 2414 -4867
rect 2444 -4867 2450 -4473
rect 2504 -4867 2510 -4473
rect 2444 -4873 2510 -4867
rect 2540 -4867 2546 -4473
rect 2600 -4867 2606 -4473
rect 2540 -4873 2606 -4867
rect 2636 -4867 2642 -4473
rect 2696 -4867 2702 -4473
rect 2636 -4873 2702 -4867
rect 2732 -4867 2738 -4473
rect 2792 -4867 2798 -4473
rect 2732 -4873 2798 -4867
rect 2828 -4867 2834 -4473
rect 2888 -4867 2894 -4473
rect 2828 -4873 2894 -4867
rect 2924 -4867 2930 -4473
rect 2984 -4867 2990 -4473
rect 2924 -4873 2990 -4867
rect 3020 -4867 3026 -4473
rect 3080 -4867 3086 -4473
rect 3020 -4873 3086 -4867
rect 3116 -4867 3122 -4473
rect 3176 -4867 3182 -4473
rect 3116 -4873 3182 -4867
rect 3212 -4867 3218 -4473
rect 3272 -4867 3278 -4473
rect 3212 -4873 3278 -4867
rect 3308 -4867 3314 -4473
rect 3368 -4867 3374 -4473
rect 3308 -4873 3374 -4867
rect 2214 -5007 2304 -4951
rect 2332 -4905 2396 -4901
rect 3314 -4905 3396 -4901
rect 2332 -4907 3396 -4905
rect 2332 -4908 3320 -4907
rect 2332 -4961 2338 -4908
rect 2390 -4961 3320 -4908
rect 2332 -4963 3320 -4961
rect 3390 -4963 3396 -4907
rect 2332 -4966 3396 -4963
rect 2332 -4967 2396 -4966
rect 3314 -4971 3396 -4966
rect 3432 -4951 3438 -4395
rect 3472 -4951 3508 -4395
rect 3432 -5007 3508 -4951
rect 2214 -5013 3508 -5007
rect 2214 -5047 2346 -5013
rect 3376 -5047 3508 -5013
rect 2214 -5083 3508 -5047
rect 2214 -5341 2356 -5083
rect 3366 -5341 3508 -5083
rect 2214 -5426 3508 -5341
rect 2214 -5551 2296 -5426
rect 2324 -5460 2409 -5454
rect 2324 -5513 2331 -5460
rect 2403 -5463 2409 -5460
rect 2403 -5513 2787 -5463
rect 2324 -5519 2787 -5513
rect 2214 -6141 2304 -5551
rect 2731 -5821 2787 -5519
rect 3312 -5776 3387 -5757
rect 3312 -5821 3322 -5776
rect 2731 -5877 3322 -5821
rect 2214 -6177 2657 -6141
rect 2214 -6211 2346 -6177
rect 2621 -6211 2657 -6177
rect 2214 -6229 2657 -6211
rect 2214 -6273 2304 -6229
rect 2731 -6263 2787 -5877
rect 3312 -5909 3322 -5877
rect 3374 -5909 3387 -5776
rect 3312 -5923 3387 -5909
rect 3418 -6141 3508 -5426
rect 3771 -5726 4056 -3290
rect 3079 -6177 3508 -6141
rect 3079 -6211 3101 -6177
rect 3376 -6211 3508 -6177
rect 3079 -6229 3508 -6211
rect 2214 -6629 2250 -6273
rect 2284 -6351 2304 -6273
rect 2492 -6319 3326 -6263
rect 3418 -6273 3508 -6229
rect 3418 -6351 3438 -6273
rect 2284 -6545 2354 -6351
rect 2408 -6545 2414 -6351
rect 2284 -6551 2414 -6545
rect 2444 -6545 2450 -6351
rect 2504 -6545 2510 -6351
rect 2444 -6551 2510 -6545
rect 2540 -6545 2546 -6351
rect 2600 -6545 2606 -6351
rect 2540 -6551 2606 -6545
rect 2636 -6545 2642 -6351
rect 2696 -6545 2702 -6351
rect 2636 -6551 2702 -6545
rect 2732 -6545 2738 -6351
rect 2792 -6545 2798 -6351
rect 2732 -6551 2798 -6545
rect 2828 -6545 2834 -6351
rect 2888 -6545 2894 -6351
rect 2828 -6551 2894 -6545
rect 2924 -6545 2930 -6351
rect 2984 -6545 2990 -6351
rect 2924 -6551 2990 -6545
rect 3020 -6545 3026 -6351
rect 3080 -6545 3086 -6351
rect 3020 -6551 3086 -6545
rect 3116 -6545 3122 -6351
rect 3176 -6545 3182 -6351
rect 3116 -6551 3182 -6545
rect 3212 -6545 3218 -6351
rect 3272 -6545 3278 -6351
rect 3212 -6551 3278 -6545
rect 3308 -6545 3314 -6351
rect 3368 -6545 3438 -6351
rect 3308 -6551 3438 -6545
rect 2284 -6629 2304 -6551
rect 2214 -6671 2304 -6629
rect 2396 -6639 3230 -6583
rect 3418 -6629 3438 -6551
rect 3472 -6629 3508 -6273
rect 2214 -6677 2798 -6671
rect 2214 -6691 2354 -6677
rect 2214 -6725 2346 -6691
rect 2214 -6755 2354 -6725
rect 2792 -6755 2798 -6677
rect 2214 -6761 2798 -6755
rect 2826 -6822 2896 -6639
rect 3418 -6671 3508 -6629
rect 2924 -6677 3508 -6671
rect 2924 -6755 2930 -6677
rect 3368 -6691 3508 -6677
rect 3376 -6725 3508 -6691
rect 3368 -6755 3508 -6725
rect 2924 -6761 3508 -6755
rect 3567 -5770 4056 -5726
rect 3567 -5909 3683 -5770
rect 3822 -5909 4056 -5770
rect 3567 -6047 4056 -5909
rect 3567 -6822 3637 -6047
rect -6172 -7150 -5411 -6864
rect 1269 -6892 3637 -6822
rect 2348 -6988 3374 -6963
rect 2348 -7150 2391 -6988
rect 3339 -7150 3374 -6988
rect -6172 -7536 -6013 -7150
rect -5627 -7536 3374 -7150
rect -6172 -7739 -5411 -7536
rect 5287 -15521 5571 -2710
rect 5974 -3009 5980 -2725
rect 6264 -3009 6270 -2725
rect 2599 -15805 5571 -15521
rect 2599 -17524 2883 -15805
rect 5980 -16163 6264 -3009
rect 3771 -16447 6264 -16163
rect 368 -17580 3619 -17524
rect 368 -17771 424 -17580
rect 606 -17656 2112 -17649
rect 606 -17685 642 -17656
rect 1967 -17685 2112 -17656
rect 606 -17719 630 -17685
rect 1980 -17719 2112 -17685
rect 606 -17729 642 -17719
rect 1967 -17729 2112 -17719
rect 606 -17735 2112 -17729
rect 368 -17827 822 -17771
rect 2022 -17781 2112 -17735
rect 368 -18898 424 -17827
rect 2022 -17868 2042 -17781
rect 498 -17874 694 -17868
rect 360 -18912 432 -18898
rect 360 -18968 368 -18912
rect 424 -18968 432 -18912
rect 360 -18974 432 -18968
rect 498 -18955 534 -17874
rect 568 -17875 694 -17874
rect 568 -18862 639 -17875
rect 692 -18862 694 -17875
rect 568 -18868 694 -18862
rect 764 -17875 822 -17868
rect 764 -18862 767 -17875
rect 820 -18862 822 -17875
rect 764 -18868 822 -18862
rect 892 -17875 950 -17868
rect 892 -18862 895 -17875
rect 948 -18862 950 -17875
rect 892 -18868 950 -18862
rect 1020 -17875 1078 -17868
rect 1020 -18862 1023 -17875
rect 1076 -18862 1078 -17875
rect 1020 -18868 1078 -18862
rect 1148 -17875 1206 -17868
rect 1148 -18862 1151 -17875
rect 1204 -18862 1206 -17875
rect 1148 -18868 1206 -18862
rect 1276 -17875 1334 -17868
rect 1276 -18862 1279 -17875
rect 1332 -18862 1334 -17875
rect 1276 -18868 1334 -18862
rect 1404 -17875 1462 -17868
rect 1404 -18862 1407 -17875
rect 1460 -18862 1462 -17875
rect 1404 -18868 1462 -18862
rect 1532 -17875 1590 -17868
rect 1532 -18862 1535 -17875
rect 1588 -18862 1590 -17875
rect 1532 -18868 1590 -18862
rect 1660 -17875 1718 -17868
rect 1660 -18862 1663 -17875
rect 1716 -18862 1718 -17875
rect 1660 -18868 1718 -18862
rect 1788 -17875 1846 -17868
rect 1788 -18862 1791 -17875
rect 1844 -18862 1846 -17875
rect 1788 -18868 1846 -18862
rect 1916 -17875 2042 -17868
rect 1916 -18862 1919 -17875
rect 1972 -18862 2042 -17875
rect 1916 -18868 2042 -18862
rect 568 -18955 578 -18868
rect 498 -19008 578 -18955
rect 614 -18909 682 -18903
rect 1904 -18907 1989 -18901
rect 1904 -18909 1911 -18907
rect 614 -18965 620 -18909
rect 676 -18965 946 -18909
rect 1896 -18960 1911 -18909
rect 1983 -18960 1989 -18907
rect 1896 -18965 1989 -18960
rect 2022 -18955 2042 -18868
rect 2076 -18955 2112 -17781
rect 614 -18971 682 -18965
rect 2022 -19008 2112 -18955
rect 498 -19017 2112 -19008
rect 498 -19051 630 -19017
rect 1980 -19051 2112 -19017
rect 498 -19087 2112 -19051
rect 498 -19341 602 -19087
rect 2008 -19341 2112 -19087
rect 498 -19377 2112 -19341
rect 498 -19411 630 -19377
rect 1980 -19411 2112 -19377
rect 498 -19427 2112 -19411
rect 498 -19473 588 -19427
rect 498 -20647 534 -19473
rect 568 -20647 588 -19473
rect 1902 -19461 1987 -19455
rect 1902 -19514 1909 -19461
rect 1981 -19514 1987 -19461
rect 1902 -19519 1987 -19514
rect 2022 -19473 2112 -19427
rect 636 -19567 694 -19560
rect 636 -20554 639 -19567
rect 692 -20554 694 -19567
rect 636 -20560 694 -20554
rect 764 -19567 822 -19560
rect 764 -20554 767 -19567
rect 820 -20554 822 -19567
rect 764 -20560 822 -20554
rect 892 -19567 950 -19560
rect 892 -20554 895 -19567
rect 948 -20554 950 -19567
rect 892 -20560 950 -20554
rect 1020 -19567 1078 -19560
rect 1020 -20554 1023 -19567
rect 1076 -20554 1078 -19567
rect 1020 -20560 1078 -20554
rect 1148 -19567 1206 -19560
rect 1148 -20554 1151 -19567
rect 1204 -20554 1206 -19567
rect 1148 -20560 1206 -20554
rect 1276 -19567 1334 -19560
rect 1276 -20554 1279 -19567
rect 1332 -20554 1334 -19567
rect 1276 -20560 1334 -20554
rect 1404 -19567 1462 -19560
rect 1404 -20554 1407 -19567
rect 1460 -20554 1462 -19567
rect 1404 -20560 1462 -20554
rect 1532 -19567 1590 -19560
rect 1532 -20554 1535 -19567
rect 1588 -20554 1590 -19567
rect 1532 -20560 1590 -20554
rect 1660 -19567 1718 -19560
rect 1660 -20554 1663 -19567
rect 1716 -20554 1718 -19567
rect 1660 -20560 1718 -20554
rect 1788 -19567 1846 -19560
rect 1788 -20554 1791 -19567
rect 1844 -20554 1846 -19567
rect 1788 -20560 1846 -20554
rect 1916 -19567 1974 -19560
rect 1916 -20554 1919 -19567
rect 1972 -20554 1974 -19567
rect 1916 -20560 1974 -20554
rect 498 -20693 588 -20647
rect 498 -20709 1227 -20693
rect 498 -20743 630 -20709
rect 1221 -20743 1227 -20709
rect 498 -20779 1227 -20743
rect 1269 -20822 1339 -20629
rect 2022 -20647 2042 -19473
rect 2076 -20647 2112 -19473
rect 2022 -20693 2112 -20647
rect 1367 -20709 2112 -20693
rect 1367 -20743 1373 -20709
rect 1980 -20743 2112 -20709
rect 1367 -20779 2112 -20743
rect 2214 -18340 2802 -18263
rect 2214 -18395 2304 -18340
rect 2834 -18385 2890 -17580
rect 3563 -17863 3619 -17580
rect 3541 -17888 3646 -17863
rect 3541 -17944 3563 -17888
rect 3619 -17944 3646 -17888
rect 3541 -17961 3646 -17944
rect 2919 -18340 3508 -18263
rect 2214 -18951 2250 -18395
rect 2284 -18951 2304 -18395
rect 2492 -18441 3326 -18385
rect 3432 -18395 3508 -18340
rect 2348 -18867 2354 -18473
rect 2408 -18867 2414 -18473
rect 2348 -18873 2414 -18867
rect 2444 -18867 2450 -18473
rect 2504 -18867 2510 -18473
rect 2444 -18873 2510 -18867
rect 2540 -18867 2546 -18473
rect 2600 -18867 2606 -18473
rect 2540 -18873 2606 -18867
rect 2636 -18867 2642 -18473
rect 2696 -18867 2702 -18473
rect 2636 -18873 2702 -18867
rect 2732 -18867 2738 -18473
rect 2792 -18867 2798 -18473
rect 2732 -18873 2798 -18867
rect 2828 -18867 2834 -18473
rect 2888 -18867 2894 -18473
rect 2828 -18873 2894 -18867
rect 2924 -18867 2930 -18473
rect 2984 -18867 2990 -18473
rect 2924 -18873 2990 -18867
rect 3020 -18867 3026 -18473
rect 3080 -18867 3086 -18473
rect 3020 -18873 3086 -18867
rect 3116 -18867 3122 -18473
rect 3176 -18867 3182 -18473
rect 3116 -18873 3182 -18867
rect 3212 -18867 3218 -18473
rect 3272 -18867 3278 -18473
rect 3212 -18873 3278 -18867
rect 3308 -18867 3314 -18473
rect 3368 -18867 3374 -18473
rect 3308 -18873 3374 -18867
rect 2214 -19007 2304 -18951
rect 2332 -18905 2396 -18901
rect 3314 -18905 3396 -18901
rect 2332 -18907 3396 -18905
rect 2332 -18908 3320 -18907
rect 2332 -18961 2338 -18908
rect 2390 -18961 3320 -18908
rect 2332 -18963 3320 -18961
rect 3390 -18963 3396 -18907
rect 2332 -18966 3396 -18963
rect 2332 -18967 2396 -18966
rect 3314 -18971 3396 -18966
rect 3432 -18951 3438 -18395
rect 3472 -18951 3508 -18395
rect 3432 -19007 3508 -18951
rect 2214 -19013 3508 -19007
rect 2214 -19047 2346 -19013
rect 3376 -19047 3508 -19013
rect 2214 -19083 3508 -19047
rect 2214 -19341 2356 -19083
rect 3366 -19341 3508 -19083
rect 2214 -19426 3508 -19341
rect 2214 -19551 2296 -19426
rect 2324 -19460 2409 -19454
rect 2324 -19513 2331 -19460
rect 2403 -19463 2409 -19460
rect 2403 -19513 2787 -19463
rect 2324 -19519 2787 -19513
rect 2214 -20141 2304 -19551
rect 2731 -19821 2787 -19519
rect 3312 -19776 3387 -19757
rect 3312 -19821 3322 -19776
rect 2731 -19877 3322 -19821
rect 2214 -20177 2657 -20141
rect 2214 -20211 2346 -20177
rect 2621 -20211 2657 -20177
rect 2214 -20229 2657 -20211
rect 2214 -20273 2304 -20229
rect 2731 -20263 2787 -19877
rect 3312 -19909 3322 -19877
rect 3374 -19909 3387 -19776
rect 3312 -19923 3387 -19909
rect 3418 -20141 3508 -19426
rect 3771 -19726 4056 -16447
rect 3079 -20177 3508 -20141
rect 3079 -20211 3101 -20177
rect 3376 -20211 3508 -20177
rect 3079 -20229 3508 -20211
rect 2214 -20629 2250 -20273
rect 2284 -20351 2304 -20273
rect 2492 -20319 3326 -20263
rect 3418 -20273 3508 -20229
rect 3418 -20351 3438 -20273
rect 2284 -20545 2354 -20351
rect 2408 -20545 2414 -20351
rect 2284 -20551 2414 -20545
rect 2444 -20545 2450 -20351
rect 2504 -20545 2510 -20351
rect 2444 -20551 2510 -20545
rect 2540 -20545 2546 -20351
rect 2600 -20545 2606 -20351
rect 2540 -20551 2606 -20545
rect 2636 -20545 2642 -20351
rect 2696 -20545 2702 -20351
rect 2636 -20551 2702 -20545
rect 2732 -20545 2738 -20351
rect 2792 -20545 2798 -20351
rect 2732 -20551 2798 -20545
rect 2828 -20545 2834 -20351
rect 2888 -20545 2894 -20351
rect 2828 -20551 2894 -20545
rect 2924 -20545 2930 -20351
rect 2984 -20545 2990 -20351
rect 2924 -20551 2990 -20545
rect 3020 -20545 3026 -20351
rect 3080 -20545 3086 -20351
rect 3020 -20551 3086 -20545
rect 3116 -20545 3122 -20351
rect 3176 -20545 3182 -20351
rect 3116 -20551 3182 -20545
rect 3212 -20545 3218 -20351
rect 3272 -20545 3278 -20351
rect 3212 -20551 3278 -20545
rect 3308 -20545 3314 -20351
rect 3368 -20545 3438 -20351
rect 3308 -20551 3438 -20545
rect 2284 -20629 2304 -20551
rect 2214 -20671 2304 -20629
rect 2396 -20639 3230 -20583
rect 3418 -20629 3438 -20551
rect 3472 -20629 3508 -20273
rect 2214 -20677 2798 -20671
rect 2214 -20691 2354 -20677
rect 2214 -20725 2346 -20691
rect 2214 -20755 2354 -20725
rect 2792 -20755 2798 -20677
rect 2214 -20761 2798 -20755
rect 2826 -20822 2896 -20639
rect 3418 -20671 3508 -20629
rect 2924 -20677 3508 -20671
rect 2924 -20755 2930 -20677
rect 3368 -20691 3508 -20677
rect 3376 -20725 3508 -20691
rect 3368 -20755 3508 -20725
rect 2924 -20761 3508 -20755
rect 3567 -19770 4056 -19726
rect 3567 -19909 3683 -19770
rect 3822 -19909 4056 -19770
rect 3567 -20047 4056 -19909
rect 3567 -20822 3637 -20047
rect -6172 -21150 -5411 -20864
rect 1269 -20892 3637 -20822
rect 2348 -20988 3374 -20963
rect 2348 -21150 2391 -20988
rect 3339 -21150 3374 -20988
rect -6172 -21536 -6013 -21150
rect -5627 -21536 3374 -21150
rect -6172 -21739 -5411 -21536
rect 7975 -29597 8259 -2710
rect 8660 -3032 8959 -3024
rect 8660 -3316 8668 -3032
rect 8952 -3316 8959 -3032
rect 8660 -3323 8959 -3316
rect 2599 -29881 8259 -29597
rect 2599 -31524 2883 -29881
rect 8668 -30327 8952 -3323
rect 3771 -30611 8952 -30327
rect 3771 -30969 4056 -30611
rect 3772 -31327 4056 -30969
rect 368 -31580 3619 -31524
rect 368 -31771 424 -31580
rect 606 -31656 2112 -31649
rect 606 -31685 642 -31656
rect 1967 -31685 2112 -31656
rect 606 -31719 630 -31685
rect 1980 -31719 2112 -31685
rect 606 -31729 642 -31719
rect 1967 -31729 2112 -31719
rect 606 -31735 2112 -31729
rect 368 -31827 822 -31771
rect 2022 -31781 2112 -31735
rect 368 -32898 424 -31827
rect 2022 -31868 2042 -31781
rect 498 -31874 694 -31868
rect 360 -32912 432 -32898
rect 360 -32968 368 -32912
rect 424 -32968 432 -32912
rect 360 -32974 432 -32968
rect 498 -32955 534 -31874
rect 568 -31875 694 -31874
rect 568 -32862 639 -31875
rect 692 -32862 694 -31875
rect 568 -32868 694 -32862
rect 764 -31875 822 -31868
rect 764 -32862 767 -31875
rect 820 -32862 822 -31875
rect 764 -32868 822 -32862
rect 892 -31875 950 -31868
rect 892 -32862 895 -31875
rect 948 -32862 950 -31875
rect 892 -32868 950 -32862
rect 1020 -31875 1078 -31868
rect 1020 -32862 1023 -31875
rect 1076 -32862 1078 -31875
rect 1020 -32868 1078 -32862
rect 1148 -31875 1206 -31868
rect 1148 -32862 1151 -31875
rect 1204 -32862 1206 -31875
rect 1148 -32868 1206 -32862
rect 1276 -31875 1334 -31868
rect 1276 -32862 1279 -31875
rect 1332 -32862 1334 -31875
rect 1276 -32868 1334 -32862
rect 1404 -31875 1462 -31868
rect 1404 -32862 1407 -31875
rect 1460 -32862 1462 -31875
rect 1404 -32868 1462 -32862
rect 1532 -31875 1590 -31868
rect 1532 -32862 1535 -31875
rect 1588 -32862 1590 -31875
rect 1532 -32868 1590 -32862
rect 1660 -31875 1718 -31868
rect 1660 -32862 1663 -31875
rect 1716 -32862 1718 -31875
rect 1660 -32868 1718 -32862
rect 1788 -31875 1846 -31868
rect 1788 -32862 1791 -31875
rect 1844 -32862 1846 -31875
rect 1788 -32868 1846 -32862
rect 1916 -31875 2042 -31868
rect 1916 -32862 1919 -31875
rect 1972 -32862 2042 -31875
rect 1916 -32868 2042 -32862
rect 568 -32955 578 -32868
rect 498 -33008 578 -32955
rect 614 -32909 682 -32903
rect 1904 -32907 1989 -32901
rect 1904 -32909 1911 -32907
rect 614 -32965 620 -32909
rect 676 -32965 946 -32909
rect 1896 -32960 1911 -32909
rect 1983 -32960 1989 -32907
rect 1896 -32965 1989 -32960
rect 2022 -32955 2042 -32868
rect 2076 -32955 2112 -31781
rect 614 -32971 682 -32965
rect 2022 -33008 2112 -32955
rect 498 -33017 2112 -33008
rect 498 -33051 630 -33017
rect 1980 -33051 2112 -33017
rect 498 -33087 2112 -33051
rect 498 -33341 602 -33087
rect 2008 -33341 2112 -33087
rect 498 -33377 2112 -33341
rect 498 -33411 630 -33377
rect 1980 -33411 2112 -33377
rect 498 -33427 2112 -33411
rect 498 -33473 588 -33427
rect 498 -34647 534 -33473
rect 568 -34647 588 -33473
rect 1902 -33461 1987 -33455
rect 1902 -33514 1909 -33461
rect 1981 -33514 1987 -33461
rect 1902 -33519 1987 -33514
rect 2022 -33473 2112 -33427
rect 636 -33567 694 -33560
rect 636 -34554 639 -33567
rect 692 -34554 694 -33567
rect 636 -34560 694 -34554
rect 764 -33567 822 -33560
rect 764 -34554 767 -33567
rect 820 -34554 822 -33567
rect 764 -34560 822 -34554
rect 892 -33567 950 -33560
rect 892 -34554 895 -33567
rect 948 -34554 950 -33567
rect 892 -34560 950 -34554
rect 1020 -33567 1078 -33560
rect 1020 -34554 1023 -33567
rect 1076 -34554 1078 -33567
rect 1020 -34560 1078 -34554
rect 1148 -33567 1206 -33560
rect 1148 -34554 1151 -33567
rect 1204 -34554 1206 -33567
rect 1148 -34560 1206 -34554
rect 1276 -33567 1334 -33560
rect 1276 -34554 1279 -33567
rect 1332 -34554 1334 -33567
rect 1276 -34560 1334 -34554
rect 1404 -33567 1462 -33560
rect 1404 -34554 1407 -33567
rect 1460 -34554 1462 -33567
rect 1404 -34560 1462 -34554
rect 1532 -33567 1590 -33560
rect 1532 -34554 1535 -33567
rect 1588 -34554 1590 -33567
rect 1532 -34560 1590 -34554
rect 1660 -33567 1718 -33560
rect 1660 -34554 1663 -33567
rect 1716 -34554 1718 -33567
rect 1660 -34560 1718 -34554
rect 1788 -33567 1846 -33560
rect 1788 -34554 1791 -33567
rect 1844 -34554 1846 -33567
rect 1788 -34560 1846 -34554
rect 1916 -33567 1974 -33560
rect 1916 -34554 1919 -33567
rect 1972 -34554 1974 -33567
rect 1916 -34560 1974 -34554
rect 498 -34693 588 -34647
rect 498 -34709 1227 -34693
rect 498 -34743 630 -34709
rect 1221 -34743 1227 -34709
rect 498 -34779 1227 -34743
rect 1269 -34822 1339 -34629
rect 2022 -34647 2042 -33473
rect 2076 -34647 2112 -33473
rect 2022 -34693 2112 -34647
rect 1367 -34709 2112 -34693
rect 1367 -34743 1373 -34709
rect 1980 -34743 2112 -34709
rect 1367 -34779 2112 -34743
rect 2214 -32340 2802 -32263
rect 2214 -32395 2304 -32340
rect 2834 -32385 2890 -31580
rect 3563 -31863 3619 -31580
rect 3541 -31888 3646 -31863
rect 3541 -31944 3563 -31888
rect 3619 -31944 3646 -31888
rect 3541 -31961 3646 -31944
rect 2919 -32340 3508 -32263
rect 2214 -32951 2250 -32395
rect 2284 -32951 2304 -32395
rect 2492 -32441 3326 -32385
rect 3432 -32395 3508 -32340
rect 2348 -32867 2354 -32473
rect 2408 -32867 2414 -32473
rect 2348 -32873 2414 -32867
rect 2444 -32867 2450 -32473
rect 2504 -32867 2510 -32473
rect 2444 -32873 2510 -32867
rect 2540 -32867 2546 -32473
rect 2600 -32867 2606 -32473
rect 2540 -32873 2606 -32867
rect 2636 -32867 2642 -32473
rect 2696 -32867 2702 -32473
rect 2636 -32873 2702 -32867
rect 2732 -32867 2738 -32473
rect 2792 -32867 2798 -32473
rect 2732 -32873 2798 -32867
rect 2828 -32867 2834 -32473
rect 2888 -32867 2894 -32473
rect 2828 -32873 2894 -32867
rect 2924 -32867 2930 -32473
rect 2984 -32867 2990 -32473
rect 2924 -32873 2990 -32867
rect 3020 -32867 3026 -32473
rect 3080 -32867 3086 -32473
rect 3020 -32873 3086 -32867
rect 3116 -32867 3122 -32473
rect 3176 -32867 3182 -32473
rect 3116 -32873 3182 -32867
rect 3212 -32867 3218 -32473
rect 3272 -32867 3278 -32473
rect 3212 -32873 3278 -32867
rect 3308 -32867 3314 -32473
rect 3368 -32867 3374 -32473
rect 3308 -32873 3374 -32867
rect 2214 -33007 2304 -32951
rect 2332 -32905 2396 -32901
rect 3314 -32905 3396 -32901
rect 2332 -32907 3396 -32905
rect 2332 -32908 3320 -32907
rect 2332 -32961 2338 -32908
rect 2390 -32961 3320 -32908
rect 2332 -32963 3320 -32961
rect 3390 -32963 3396 -32907
rect 2332 -32966 3396 -32963
rect 2332 -32967 2396 -32966
rect 3314 -32971 3396 -32966
rect 3432 -32951 3438 -32395
rect 3472 -32951 3508 -32395
rect 3432 -33007 3508 -32951
rect 2214 -33013 3508 -33007
rect 2214 -33047 2346 -33013
rect 3376 -33047 3508 -33013
rect 2214 -33083 3508 -33047
rect 2214 -33341 2356 -33083
rect 3366 -33341 3508 -33083
rect 2214 -33426 3508 -33341
rect 2214 -33551 2296 -33426
rect 2324 -33460 2409 -33454
rect 2324 -33513 2331 -33460
rect 2403 -33463 2409 -33460
rect 2403 -33513 2787 -33463
rect 2324 -33519 2787 -33513
rect 2214 -34141 2304 -33551
rect 2731 -33821 2787 -33519
rect 3312 -33776 3387 -33757
rect 3312 -33821 3322 -33776
rect 2731 -33877 3322 -33821
rect 2214 -34177 2657 -34141
rect 2214 -34211 2346 -34177
rect 2621 -34211 2657 -34177
rect 2214 -34229 2657 -34211
rect 2214 -34273 2304 -34229
rect 2731 -34263 2787 -33877
rect 3312 -33909 3322 -33877
rect 3374 -33909 3387 -33776
rect 3312 -33923 3387 -33909
rect 3418 -34141 3508 -33426
rect 3771 -33726 4056 -31327
rect 3079 -34177 3508 -34141
rect 3079 -34211 3101 -34177
rect 3376 -34211 3508 -34177
rect 3079 -34229 3508 -34211
rect 2214 -34629 2250 -34273
rect 2284 -34351 2304 -34273
rect 2492 -34319 3326 -34263
rect 3418 -34273 3508 -34229
rect 3418 -34351 3438 -34273
rect 2284 -34545 2354 -34351
rect 2408 -34545 2414 -34351
rect 2284 -34551 2414 -34545
rect 2444 -34545 2450 -34351
rect 2504 -34545 2510 -34351
rect 2444 -34551 2510 -34545
rect 2540 -34545 2546 -34351
rect 2600 -34545 2606 -34351
rect 2540 -34551 2606 -34545
rect 2636 -34545 2642 -34351
rect 2696 -34545 2702 -34351
rect 2636 -34551 2702 -34545
rect 2732 -34545 2738 -34351
rect 2792 -34545 2798 -34351
rect 2732 -34551 2798 -34545
rect 2828 -34545 2834 -34351
rect 2888 -34545 2894 -34351
rect 2828 -34551 2894 -34545
rect 2924 -34545 2930 -34351
rect 2984 -34545 2990 -34351
rect 2924 -34551 2990 -34545
rect 3020 -34545 3026 -34351
rect 3080 -34545 3086 -34351
rect 3020 -34551 3086 -34545
rect 3116 -34545 3122 -34351
rect 3176 -34545 3182 -34351
rect 3116 -34551 3182 -34545
rect 3212 -34545 3218 -34351
rect 3272 -34545 3278 -34351
rect 3212 -34551 3278 -34545
rect 3308 -34545 3314 -34351
rect 3368 -34545 3438 -34351
rect 3308 -34551 3438 -34545
rect 2284 -34629 2304 -34551
rect 2214 -34671 2304 -34629
rect 2396 -34639 3230 -34583
rect 3418 -34629 3438 -34551
rect 3472 -34629 3508 -34273
rect 2214 -34677 2798 -34671
rect 2214 -34691 2354 -34677
rect 2214 -34725 2346 -34691
rect 2214 -34755 2354 -34725
rect 2792 -34755 2798 -34677
rect 2214 -34761 2798 -34755
rect 2826 -34822 2896 -34639
rect 3418 -34671 3508 -34629
rect 2924 -34677 3508 -34671
rect 2924 -34755 2930 -34677
rect 3368 -34691 3508 -34677
rect 3376 -34725 3508 -34691
rect 3368 -34755 3508 -34725
rect 2924 -34761 3508 -34755
rect 3567 -33770 4056 -33726
rect 3567 -33909 3683 -33770
rect 3822 -33909 4056 -33770
rect 3567 -34047 4056 -33909
rect 3567 -34822 3637 -34047
rect -6172 -35150 -5411 -34864
rect 1269 -34892 3637 -34822
rect 2348 -34988 3374 -34963
rect 2348 -35150 2391 -34988
rect 3339 -35150 3374 -34988
rect -6172 -35536 -6013 -35150
rect -5627 -35536 3374 -35150
rect -6172 -35739 -5411 -35536
rect 10663 -42890 10947 -2710
rect 11384 -2712 11474 -2670
rect 12820 -2670 12840 -2532
rect 12874 -2670 12950 -2532
rect 12984 -2670 13004 -2532
rect 14350 -2532 14440 -2490
rect 13080 -2572 13512 -2566
rect 13080 -2630 13088 -2572
rect 13504 -2630 13512 -2572
rect 13080 -2636 13512 -2630
rect 13842 -2572 14274 -2566
rect 13842 -2630 13850 -2572
rect 14266 -2630 14274 -2572
rect 13842 -2636 14274 -2630
rect 12820 -2712 13004 -2670
rect 14350 -2670 14370 -2532
rect 14404 -2670 14440 -2532
rect 14350 -2712 14440 -2670
rect 11384 -2732 14440 -2712
rect 11384 -2766 11516 -2732
rect 12778 -2766 13046 -2732
rect 14308 -2766 14440 -2732
rect 11384 -2802 14440 -2766
rect 11350 -3476 11356 -3192
rect 11640 -3476 11646 -3192
rect 2599 -43174 10947 -42890
rect 2599 -45524 2883 -43174
rect 11356 -43796 11640 -3476
rect 41396 -11731 41568 489
rect 40960 -11743 42222 -11731
rect 40960 -11777 41068 -11743
rect 42114 -11777 42222 -11743
rect 40960 -11789 42222 -11777
rect 40960 -11839 41018 -11789
rect 40960 -24589 40972 -11839
rect 41006 -24589 41018 -11839
rect 42032 -11849 42133 -11830
rect 41191 -11867 41991 -11859
rect 41191 -11921 41203 -11867
rect 41979 -11921 41991 -11867
rect 41094 -11957 41150 -11923
rect 41191 -11929 41991 -11921
rect 42032 -11916 42050 -11849
rect 42114 -11916 42133 -11849
rect 42032 -11934 42133 -11916
rect 42164 -11839 42222 -11789
rect 42032 -11957 42088 -11934
rect 41094 -11989 42088 -11957
rect 41094 -12115 41150 -11989
rect 41191 -12025 41991 -12017
rect 41191 -12079 41203 -12025
rect 41979 -12079 41991 -12025
rect 41191 -12087 41991 -12079
rect 42032 -12115 42088 -11989
rect 41094 -12147 42088 -12115
rect 41094 -12273 41150 -12147
rect 41191 -12183 41991 -12175
rect 41191 -12237 41203 -12183
rect 41979 -12237 41991 -12183
rect 41191 -12245 41991 -12237
rect 42032 -12273 42088 -12147
rect 41094 -12305 42088 -12273
rect 41094 -12431 41150 -12305
rect 41191 -12341 41991 -12333
rect 41191 -12395 41203 -12341
rect 41979 -12395 41991 -12341
rect 41191 -12403 41991 -12395
rect 42032 -12431 42088 -12305
rect 41094 -12463 42088 -12431
rect 41094 -12589 41150 -12463
rect 41191 -12499 41991 -12491
rect 41191 -12553 41203 -12499
rect 41979 -12553 41991 -12499
rect 41191 -12561 41991 -12553
rect 42032 -12589 42088 -12463
rect 41094 -12621 42088 -12589
rect 41094 -12747 41150 -12621
rect 41191 -12657 41991 -12649
rect 41191 -12711 41203 -12657
rect 41979 -12711 41991 -12657
rect 41191 -12719 41991 -12711
rect 42032 -12747 42088 -12621
rect 41094 -12779 42088 -12747
rect 41094 -12905 41150 -12779
rect 41191 -12815 41991 -12807
rect 41191 -12869 41203 -12815
rect 41979 -12869 41991 -12815
rect 41191 -12877 41991 -12869
rect 42032 -12905 42088 -12779
rect 41094 -12937 42088 -12905
rect 41094 -13063 41150 -12937
rect 41191 -12973 41991 -12965
rect 41191 -13027 41203 -12973
rect 41979 -13027 41991 -12973
rect 41191 -13035 41991 -13027
rect 42032 -13063 42088 -12937
rect 41094 -13095 42088 -13063
rect 41094 -13221 41150 -13095
rect 41191 -13131 41991 -13123
rect 41191 -13185 41203 -13131
rect 41979 -13185 41991 -13131
rect 41191 -13193 41991 -13185
rect 42032 -13221 42088 -13095
rect 41094 -13253 42088 -13221
rect 41094 -13379 41150 -13253
rect 41191 -13289 41991 -13281
rect 41191 -13343 41203 -13289
rect 41979 -13343 41991 -13289
rect 41191 -13351 41991 -13343
rect 42032 -13379 42088 -13253
rect 41094 -13411 42088 -13379
rect 41094 -13537 41150 -13411
rect 41191 -13447 41991 -13439
rect 41191 -13501 41203 -13447
rect 41979 -13501 41991 -13447
rect 41191 -13509 41991 -13501
rect 42032 -13537 42088 -13411
rect 41094 -13569 42088 -13537
rect 41094 -13695 41150 -13569
rect 41191 -13605 41991 -13597
rect 41191 -13659 41203 -13605
rect 41979 -13659 41991 -13605
rect 41191 -13667 41991 -13659
rect 42032 -13695 42088 -13569
rect 41094 -13727 42088 -13695
rect 41094 -13853 41150 -13727
rect 41191 -13763 41991 -13755
rect 41191 -13817 41203 -13763
rect 41979 -13817 41991 -13763
rect 41191 -13825 41991 -13817
rect 42032 -13853 42088 -13727
rect 41094 -13885 42088 -13853
rect 41094 -14011 41150 -13885
rect 41191 -13921 41991 -13913
rect 41191 -13975 41203 -13921
rect 41979 -13975 41991 -13921
rect 41191 -13983 41991 -13975
rect 42032 -14011 42088 -13885
rect 41094 -14043 42088 -14011
rect 41094 -14169 41150 -14043
rect 41191 -14079 41991 -14071
rect 41191 -14133 41203 -14079
rect 41979 -14133 41991 -14079
rect 41191 -14141 41991 -14133
rect 42032 -14169 42088 -14043
rect 41094 -14201 42088 -14169
rect 41094 -14327 41150 -14201
rect 41191 -14237 41991 -14229
rect 41191 -14291 41203 -14237
rect 41979 -14291 41991 -14237
rect 41191 -14299 41991 -14291
rect 42032 -14327 42088 -14201
rect 41094 -14359 42088 -14327
rect 41094 -14485 41150 -14359
rect 41191 -14395 41991 -14387
rect 41191 -14449 41203 -14395
rect 41979 -14449 41991 -14395
rect 41191 -14457 41991 -14449
rect 42032 -14485 42088 -14359
rect 41094 -14517 42088 -14485
rect 41094 -14643 41150 -14517
rect 41191 -14553 41991 -14545
rect 41191 -14607 41203 -14553
rect 41979 -14607 41991 -14553
rect 41191 -14615 41991 -14607
rect 42032 -14643 42088 -14517
rect 41094 -14675 42088 -14643
rect 41094 -14801 41150 -14675
rect 41191 -14711 41991 -14703
rect 41191 -14765 41203 -14711
rect 41979 -14765 41991 -14711
rect 41191 -14773 41991 -14765
rect 42032 -14801 42088 -14675
rect 41094 -14833 42088 -14801
rect 41094 -14959 41150 -14833
rect 41191 -14869 41991 -14861
rect 41191 -14923 41203 -14869
rect 41979 -14923 41991 -14869
rect 41191 -14931 41991 -14923
rect 42032 -14959 42088 -14833
rect 41094 -14991 42088 -14959
rect 41094 -15117 41150 -14991
rect 41191 -15027 41991 -15019
rect 41191 -15081 41203 -15027
rect 41979 -15081 41991 -15027
rect 41191 -15089 41991 -15081
rect 42032 -15117 42088 -14991
rect 41094 -15149 42088 -15117
rect 41094 -15275 41150 -15149
rect 41191 -15185 41991 -15177
rect 41191 -15239 41203 -15185
rect 41979 -15239 41991 -15185
rect 41191 -15247 41991 -15239
rect 42032 -15275 42088 -15149
rect 41094 -15307 42088 -15275
rect 41094 -15433 41150 -15307
rect 41191 -15343 41991 -15335
rect 41191 -15397 41203 -15343
rect 41979 -15397 41991 -15343
rect 41191 -15405 41991 -15397
rect 42032 -15433 42088 -15307
rect 41094 -15465 42088 -15433
rect 41094 -15591 41150 -15465
rect 41191 -15501 41991 -15493
rect 41191 -15555 41203 -15501
rect 41979 -15555 41991 -15501
rect 41191 -15563 41991 -15555
rect 42032 -15591 42088 -15465
rect 41094 -15623 42088 -15591
rect 41094 -15749 41150 -15623
rect 41191 -15659 41991 -15651
rect 41191 -15713 41203 -15659
rect 41979 -15713 41991 -15659
rect 41191 -15721 41991 -15713
rect 42032 -15749 42088 -15623
rect 41094 -15781 42088 -15749
rect 41094 -15907 41150 -15781
rect 41191 -15817 41991 -15809
rect 41191 -15871 41203 -15817
rect 41979 -15871 41991 -15817
rect 41191 -15879 41991 -15871
rect 42032 -15907 42088 -15781
rect 41094 -15939 42088 -15907
rect 41094 -16065 41150 -15939
rect 41191 -15975 41991 -15967
rect 41191 -16029 41203 -15975
rect 41979 -16029 41991 -15975
rect 41191 -16037 41991 -16029
rect 42032 -16065 42088 -15939
rect 41094 -16097 42088 -16065
rect 41094 -16223 41150 -16097
rect 41191 -16133 41991 -16125
rect 41191 -16187 41203 -16133
rect 41979 -16187 41991 -16133
rect 41191 -16195 41991 -16187
rect 42032 -16223 42088 -16097
rect 41094 -16255 42088 -16223
rect 41094 -16381 41150 -16255
rect 41191 -16291 41991 -16283
rect 41191 -16345 41203 -16291
rect 41979 -16345 41991 -16291
rect 41191 -16353 41991 -16345
rect 42032 -16381 42088 -16255
rect 41094 -16413 42088 -16381
rect 41094 -16539 41150 -16413
rect 41191 -16449 41991 -16441
rect 41191 -16503 41203 -16449
rect 41979 -16503 41991 -16449
rect 41191 -16511 41991 -16503
rect 42032 -16539 42088 -16413
rect 41094 -16571 42088 -16539
rect 41094 -16697 41150 -16571
rect 41191 -16607 41991 -16599
rect 41191 -16661 41203 -16607
rect 41979 -16661 41991 -16607
rect 41191 -16669 41991 -16661
rect 42032 -16697 42088 -16571
rect 41094 -16729 42088 -16697
rect 41094 -16855 41150 -16729
rect 41191 -16765 41991 -16757
rect 41191 -16819 41203 -16765
rect 41979 -16819 41991 -16765
rect 41191 -16827 41991 -16819
rect 42032 -16855 42088 -16729
rect 41094 -16887 42088 -16855
rect 41094 -17013 41150 -16887
rect 41191 -16923 41991 -16915
rect 41191 -16977 41203 -16923
rect 41979 -16977 41991 -16923
rect 41191 -16985 41991 -16977
rect 42032 -17013 42088 -16887
rect 41094 -17045 42088 -17013
rect 41094 -17171 41150 -17045
rect 41191 -17081 41991 -17073
rect 41191 -17135 41203 -17081
rect 41979 -17135 41991 -17081
rect 41191 -17143 41991 -17135
rect 42032 -17171 42088 -17045
rect 41094 -17203 42088 -17171
rect 41094 -17329 41150 -17203
rect 41191 -17239 41991 -17231
rect 41191 -17293 41203 -17239
rect 41979 -17293 41991 -17239
rect 41191 -17301 41991 -17293
rect 42032 -17329 42088 -17203
rect 41094 -17361 42088 -17329
rect 41094 -17487 41150 -17361
rect 41191 -17397 41991 -17389
rect 41191 -17451 41203 -17397
rect 41979 -17451 41991 -17397
rect 41191 -17459 41991 -17451
rect 42032 -17487 42088 -17361
rect 41094 -17519 42088 -17487
rect 41094 -17645 41150 -17519
rect 41191 -17555 41991 -17547
rect 41191 -17609 41203 -17555
rect 41979 -17609 41991 -17555
rect 41191 -17617 41991 -17609
rect 42032 -17645 42088 -17519
rect 41094 -17677 42088 -17645
rect 41094 -17803 41150 -17677
rect 41191 -17713 41991 -17705
rect 41191 -17767 41203 -17713
rect 41979 -17767 41991 -17713
rect 41191 -17775 41991 -17767
rect 42032 -17803 42088 -17677
rect 41094 -17835 42088 -17803
rect 41094 -17961 41150 -17835
rect 41191 -17871 41991 -17863
rect 41191 -17925 41203 -17871
rect 41979 -17925 41991 -17871
rect 41191 -17933 41991 -17925
rect 42032 -17961 42088 -17835
rect 41094 -17993 42088 -17961
rect 41094 -18119 41150 -17993
rect 41191 -18029 41991 -18021
rect 41191 -18083 41203 -18029
rect 41979 -18083 41991 -18029
rect 41191 -18091 41991 -18083
rect 42032 -18119 42088 -17993
rect 41094 -18151 42088 -18119
rect 41094 -18277 41150 -18151
rect 41191 -18187 41991 -18179
rect 41191 -18241 41203 -18187
rect 41979 -18241 41991 -18187
rect 41191 -18249 41991 -18241
rect 42032 -18277 42088 -18151
rect 41094 -18309 42088 -18277
rect 41094 -18435 41150 -18309
rect 41191 -18345 41991 -18337
rect 41191 -18399 41203 -18345
rect 41979 -18399 41991 -18345
rect 41191 -18407 41991 -18399
rect 42032 -18435 42088 -18309
rect 41094 -18467 42088 -18435
rect 41094 -18593 41150 -18467
rect 41191 -18503 41991 -18495
rect 41191 -18557 41203 -18503
rect 41979 -18557 41991 -18503
rect 41191 -18565 41991 -18557
rect 42032 -18593 42088 -18467
rect 41094 -18625 42088 -18593
rect 41094 -18751 41150 -18625
rect 41191 -18661 41991 -18653
rect 41191 -18715 41203 -18661
rect 41979 -18715 41991 -18661
rect 41191 -18723 41991 -18715
rect 42032 -18751 42088 -18625
rect 41094 -18783 42088 -18751
rect 41094 -18909 41150 -18783
rect 41191 -18819 41991 -18811
rect 41191 -18873 41203 -18819
rect 41979 -18873 41991 -18819
rect 41191 -18881 41991 -18873
rect 42032 -18909 42088 -18783
rect 41094 -18941 42088 -18909
rect 41094 -19067 41150 -18941
rect 41191 -18977 41991 -18969
rect 41191 -19031 41203 -18977
rect 41979 -19031 41991 -18977
rect 41191 -19039 41991 -19031
rect 42032 -19067 42088 -18941
rect 41094 -19099 42088 -19067
rect 41094 -19225 41150 -19099
rect 41191 -19135 41991 -19127
rect 41191 -19189 41203 -19135
rect 41979 -19189 41991 -19135
rect 41191 -19197 41991 -19189
rect 42032 -19225 42088 -19099
rect 41094 -19257 42088 -19225
rect 41094 -19383 41150 -19257
rect 41191 -19293 41991 -19285
rect 41191 -19347 41203 -19293
rect 41979 -19347 41991 -19293
rect 41191 -19355 41991 -19347
rect 42032 -19383 42088 -19257
rect 41094 -19415 42088 -19383
rect 41094 -19541 41150 -19415
rect 41191 -19451 41991 -19443
rect 41191 -19505 41203 -19451
rect 41979 -19505 41991 -19451
rect 41191 -19513 41991 -19505
rect 42032 -19541 42088 -19415
rect 41094 -19573 42088 -19541
rect 41094 -19699 41150 -19573
rect 41191 -19609 41991 -19601
rect 41191 -19663 41203 -19609
rect 41979 -19663 41991 -19609
rect 41191 -19671 41991 -19663
rect 42032 -19699 42088 -19573
rect 41094 -19731 42088 -19699
rect 41094 -19857 41150 -19731
rect 41191 -19767 41991 -19759
rect 41191 -19821 41203 -19767
rect 41979 -19821 41991 -19767
rect 41191 -19829 41991 -19821
rect 42032 -19857 42088 -19731
rect 41094 -19889 42088 -19857
rect 41094 -20015 41150 -19889
rect 41191 -19925 41991 -19917
rect 41191 -19979 41203 -19925
rect 41979 -19979 41991 -19925
rect 41191 -19987 41991 -19979
rect 42032 -20015 42088 -19889
rect 41094 -20047 42088 -20015
rect 41094 -20173 41150 -20047
rect 41191 -20083 41991 -20075
rect 41191 -20137 41203 -20083
rect 41979 -20137 41991 -20083
rect 41191 -20145 41991 -20137
rect 42032 -20173 42088 -20047
rect 41094 -20205 42088 -20173
rect 41094 -20331 41150 -20205
rect 41191 -20241 41991 -20233
rect 41191 -20295 41203 -20241
rect 41979 -20295 41991 -20241
rect 41191 -20303 41991 -20295
rect 42032 -20331 42088 -20205
rect 41094 -20363 42088 -20331
rect 41094 -20489 41150 -20363
rect 41191 -20399 41991 -20391
rect 41191 -20453 41203 -20399
rect 41979 -20453 41991 -20399
rect 41191 -20461 41991 -20453
rect 42032 -20489 42088 -20363
rect 41094 -20521 42088 -20489
rect 41094 -20647 41150 -20521
rect 41191 -20557 41991 -20549
rect 41191 -20611 41203 -20557
rect 41979 -20611 41991 -20557
rect 41191 -20619 41991 -20611
rect 42032 -20647 42088 -20521
rect 41094 -20679 42088 -20647
rect 41094 -20805 41150 -20679
rect 41191 -20715 41991 -20707
rect 41191 -20769 41203 -20715
rect 41979 -20769 41991 -20715
rect 41191 -20777 41991 -20769
rect 42032 -20805 42088 -20679
rect 41094 -20837 42088 -20805
rect 41094 -20963 41150 -20837
rect 41191 -20873 41991 -20865
rect 41191 -20927 41203 -20873
rect 41979 -20927 41991 -20873
rect 41191 -20935 41991 -20927
rect 42032 -20963 42088 -20837
rect 41094 -20995 42088 -20963
rect 41094 -21121 41150 -20995
rect 41191 -21031 41991 -21023
rect 41191 -21085 41203 -21031
rect 41979 -21085 41991 -21031
rect 41191 -21093 41991 -21085
rect 42032 -21121 42088 -20995
rect 41094 -21153 42088 -21121
rect 41094 -21279 41150 -21153
rect 41191 -21189 41991 -21181
rect 41191 -21243 41203 -21189
rect 41979 -21243 41991 -21189
rect 41191 -21251 41991 -21243
rect 42032 -21279 42088 -21153
rect 41094 -21311 42088 -21279
rect 41094 -21437 41150 -21311
rect 41191 -21347 41991 -21339
rect 41191 -21401 41203 -21347
rect 41979 -21401 41991 -21347
rect 41191 -21409 41991 -21401
rect 42032 -21437 42088 -21311
rect 41094 -21469 42088 -21437
rect 41094 -21595 41150 -21469
rect 41191 -21505 41991 -21497
rect 41191 -21559 41203 -21505
rect 41979 -21559 41991 -21505
rect 41191 -21567 41991 -21559
rect 42032 -21595 42088 -21469
rect 41094 -21627 42088 -21595
rect 41094 -21753 41150 -21627
rect 41191 -21663 41991 -21655
rect 41191 -21717 41203 -21663
rect 41979 -21717 41991 -21663
rect 41191 -21725 41991 -21717
rect 42032 -21753 42088 -21627
rect 41094 -21785 42088 -21753
rect 41094 -21911 41150 -21785
rect 41191 -21821 41991 -21813
rect 41191 -21875 41203 -21821
rect 41979 -21875 41991 -21821
rect 41191 -21883 41991 -21875
rect 42032 -21911 42088 -21785
rect 41094 -21943 42088 -21911
rect 41094 -22069 41150 -21943
rect 41191 -21979 41991 -21971
rect 41191 -22033 41203 -21979
rect 41979 -22033 41991 -21979
rect 41191 -22041 41991 -22033
rect 42032 -22069 42088 -21943
rect 41094 -22101 42088 -22069
rect 41094 -22227 41150 -22101
rect 41191 -22137 41991 -22129
rect 41191 -22191 41203 -22137
rect 41979 -22191 41991 -22137
rect 41191 -22199 41991 -22191
rect 42032 -22227 42088 -22101
rect 41094 -22259 42088 -22227
rect 41094 -22385 41150 -22259
rect 41191 -22295 41991 -22287
rect 41191 -22349 41203 -22295
rect 41979 -22349 41991 -22295
rect 41191 -22357 41991 -22349
rect 42032 -22385 42088 -22259
rect 41094 -22417 42088 -22385
rect 41094 -22543 41150 -22417
rect 41191 -22453 41991 -22445
rect 41191 -22507 41203 -22453
rect 41979 -22507 41991 -22453
rect 41191 -22515 41991 -22507
rect 42032 -22543 42088 -22417
rect 41094 -22575 42088 -22543
rect 41094 -22701 41150 -22575
rect 41191 -22611 41991 -22603
rect 41191 -22665 41203 -22611
rect 41979 -22665 41991 -22611
rect 41191 -22673 41991 -22665
rect 42032 -22701 42088 -22575
rect 41094 -22733 42088 -22701
rect 41094 -22859 41150 -22733
rect 41191 -22769 41991 -22761
rect 41191 -22823 41203 -22769
rect 41979 -22823 41991 -22769
rect 41191 -22831 41991 -22823
rect 42032 -22859 42088 -22733
rect 41094 -22891 42088 -22859
rect 41094 -23017 41150 -22891
rect 41191 -22927 41991 -22919
rect 41191 -22981 41203 -22927
rect 41979 -22981 41991 -22927
rect 41191 -22989 41991 -22981
rect 42032 -23017 42088 -22891
rect 41094 -23049 42088 -23017
rect 41094 -23175 41150 -23049
rect 41191 -23085 41991 -23077
rect 41191 -23139 41203 -23085
rect 41979 -23139 41991 -23085
rect 41191 -23147 41991 -23139
rect 42032 -23175 42088 -23049
rect 41094 -23207 42088 -23175
rect 41094 -23333 41150 -23207
rect 41191 -23243 41991 -23235
rect 41191 -23297 41203 -23243
rect 41979 -23297 41991 -23243
rect 41191 -23305 41991 -23297
rect 42032 -23333 42088 -23207
rect 41094 -23365 42088 -23333
rect 41094 -23491 41150 -23365
rect 41191 -23401 41991 -23393
rect 41191 -23455 41203 -23401
rect 41979 -23455 41991 -23401
rect 41191 -23463 41991 -23455
rect 42032 -23491 42088 -23365
rect 41094 -23523 42088 -23491
rect 41094 -23649 41150 -23523
rect 41191 -23559 41991 -23551
rect 41191 -23613 41203 -23559
rect 41979 -23613 41991 -23559
rect 41191 -23621 41991 -23613
rect 42032 -23649 42088 -23523
rect 41094 -23681 42088 -23649
rect 41094 -23807 41150 -23681
rect 41191 -23717 41991 -23709
rect 41191 -23771 41203 -23717
rect 41979 -23771 41991 -23717
rect 41191 -23779 41991 -23771
rect 42032 -23807 42088 -23681
rect 41094 -23839 42088 -23807
rect 41094 -23965 41150 -23839
rect 41191 -23875 41991 -23867
rect 41191 -23929 41203 -23875
rect 41979 -23929 41991 -23875
rect 41191 -23937 41991 -23929
rect 42032 -23965 42088 -23839
rect 41094 -23997 42088 -23965
rect 41094 -24123 41150 -23997
rect 41191 -24033 41991 -24025
rect 41191 -24087 41203 -24033
rect 41979 -24087 41991 -24033
rect 41191 -24095 41991 -24087
rect 42032 -24123 42088 -23997
rect 41094 -24155 42088 -24123
rect 41094 -24281 41150 -24155
rect 41191 -24191 41991 -24183
rect 41191 -24245 41203 -24191
rect 41979 -24245 41991 -24191
rect 41191 -24253 41991 -24245
rect 42032 -24281 42088 -24155
rect 41094 -24313 42088 -24281
rect 41094 -24439 41150 -24313
rect 41191 -24349 41991 -24341
rect 41191 -24403 41203 -24349
rect 41979 -24403 41991 -24349
rect 41191 -24411 41991 -24403
rect 42032 -24439 42088 -24313
rect 41094 -24471 42088 -24439
rect 41094 -24505 41150 -24471
rect 41191 -24507 41991 -24499
rect 42032 -24505 42088 -24471
rect 41191 -24561 41203 -24507
rect 41979 -24561 41991 -24507
rect 41191 -24569 41991 -24561
rect 40960 -24639 41018 -24589
rect 42164 -24589 42176 -11839
rect 42210 -24589 42222 -11839
rect 42164 -24639 42222 -24589
rect 40960 -24651 42222 -24639
rect 40960 -24685 41068 -24651
rect 42114 -24685 42222 -24651
rect 40960 -24697 42222 -24685
rect 40952 -25834 42196 -25776
rect 40952 -38684 41010 -25834
rect 41174 -25912 41974 -25905
rect 41174 -25966 41186 -25912
rect 41962 -25966 41974 -25912
rect 41086 -26047 41142 -25968
rect 41174 -25973 41974 -25966
rect 42006 -25946 42105 -25938
rect 41042 -26056 41142 -26047
rect 41042 -26151 41053 -26056
rect 41128 -26151 41142 -26056
rect 42006 -26014 42014 -25946
rect 42098 -26014 42105 -25946
rect 42006 -26023 42105 -26014
rect 41174 -26070 41974 -26063
rect 41174 -26124 41186 -26070
rect 41962 -26124 41974 -26070
rect 41174 -26131 41974 -26124
rect 41042 -26159 41142 -26151
rect 41086 -38550 41142 -26159
rect 41174 -26228 41974 -26221
rect 41174 -26282 41186 -26228
rect 41962 -26282 41974 -26228
rect 41174 -26289 41974 -26282
rect 41174 -26386 41974 -26379
rect 41174 -26440 41186 -26386
rect 41962 -26440 41974 -26386
rect 41174 -26447 41974 -26440
rect 41174 -26544 41974 -26537
rect 41174 -26598 41186 -26544
rect 41962 -26598 41974 -26544
rect 41174 -26605 41974 -26598
rect 41174 -26702 41974 -26695
rect 41174 -26756 41186 -26702
rect 41962 -26756 41974 -26702
rect 41174 -26763 41974 -26756
rect 41174 -26860 41974 -26853
rect 41174 -26914 41186 -26860
rect 41962 -26914 41974 -26860
rect 41174 -26921 41974 -26914
rect 41174 -27018 41974 -27011
rect 41174 -27072 41186 -27018
rect 41962 -27072 41974 -27018
rect 41174 -27079 41974 -27072
rect 41174 -27176 41974 -27169
rect 41174 -27230 41186 -27176
rect 41962 -27230 41974 -27176
rect 41174 -27237 41974 -27230
rect 41174 -27334 41974 -27327
rect 41174 -27388 41186 -27334
rect 41962 -27388 41974 -27334
rect 41174 -27395 41974 -27388
rect 41174 -27492 41974 -27485
rect 41174 -27546 41186 -27492
rect 41962 -27546 41974 -27492
rect 41174 -27553 41974 -27546
rect 41174 -27650 41974 -27643
rect 41174 -27704 41186 -27650
rect 41962 -27704 41974 -27650
rect 41174 -27711 41974 -27704
rect 41174 -27808 41974 -27801
rect 41174 -27862 41186 -27808
rect 41962 -27862 41974 -27808
rect 41174 -27869 41974 -27862
rect 41174 -27966 41974 -27959
rect 41174 -28020 41186 -27966
rect 41962 -28020 41974 -27966
rect 41174 -28027 41974 -28020
rect 41174 -28124 41974 -28117
rect 41174 -28178 41186 -28124
rect 41962 -28178 41974 -28124
rect 41174 -28185 41974 -28178
rect 41174 -28282 41974 -28275
rect 41174 -28336 41186 -28282
rect 41962 -28336 41974 -28282
rect 41174 -28343 41974 -28336
rect 41174 -28440 41974 -28433
rect 41174 -28494 41186 -28440
rect 41962 -28494 41974 -28440
rect 41174 -28501 41974 -28494
rect 41174 -28598 41974 -28591
rect 41174 -28652 41186 -28598
rect 41962 -28652 41974 -28598
rect 41174 -28659 41974 -28652
rect 41174 -28756 41974 -28749
rect 41174 -28810 41186 -28756
rect 41962 -28810 41974 -28756
rect 41174 -28817 41974 -28810
rect 41174 -28914 41974 -28907
rect 41174 -28968 41186 -28914
rect 41962 -28968 41974 -28914
rect 41174 -28975 41974 -28968
rect 41174 -29072 41974 -29065
rect 41174 -29126 41186 -29072
rect 41962 -29126 41974 -29072
rect 41174 -29133 41974 -29126
rect 41174 -29230 41974 -29223
rect 41174 -29284 41186 -29230
rect 41962 -29284 41974 -29230
rect 41174 -29291 41974 -29284
rect 41174 -29388 41974 -29381
rect 41174 -29442 41186 -29388
rect 41962 -29442 41974 -29388
rect 41174 -29449 41974 -29442
rect 41174 -29546 41974 -29539
rect 41174 -29600 41186 -29546
rect 41962 -29600 41974 -29546
rect 41174 -29607 41974 -29600
rect 41174 -29704 41974 -29697
rect 41174 -29758 41186 -29704
rect 41962 -29758 41974 -29704
rect 41174 -29765 41974 -29758
rect 41174 -29862 41974 -29855
rect 41174 -29916 41186 -29862
rect 41962 -29916 41974 -29862
rect 41174 -29923 41974 -29916
rect 41174 -30020 41974 -30013
rect 41174 -30074 41186 -30020
rect 41962 -30074 41974 -30020
rect 41174 -30081 41974 -30074
rect 41174 -30178 41974 -30171
rect 41174 -30232 41186 -30178
rect 41962 -30232 41974 -30178
rect 41174 -30239 41974 -30232
rect 41174 -30336 41974 -30329
rect 41174 -30390 41186 -30336
rect 41962 -30390 41974 -30336
rect 41174 -30397 41974 -30390
rect 41174 -30494 41974 -30487
rect 41174 -30548 41186 -30494
rect 41962 -30548 41974 -30494
rect 41174 -30555 41974 -30548
rect 41174 -30652 41974 -30645
rect 41174 -30706 41186 -30652
rect 41962 -30706 41974 -30652
rect 41174 -30713 41974 -30706
rect 41174 -30810 41974 -30803
rect 41174 -30864 41186 -30810
rect 41962 -30864 41974 -30810
rect 41174 -30871 41974 -30864
rect 41174 -30968 41974 -30961
rect 41174 -31022 41186 -30968
rect 41962 -31022 41974 -30968
rect 41174 -31029 41974 -31022
rect 41174 -31126 41974 -31119
rect 41174 -31180 41186 -31126
rect 41962 -31180 41974 -31126
rect 41174 -31187 41974 -31180
rect 41174 -31284 41974 -31277
rect 41174 -31338 41186 -31284
rect 41962 -31338 41974 -31284
rect 41174 -31345 41974 -31338
rect 41174 -31442 41974 -31435
rect 41174 -31496 41186 -31442
rect 41962 -31496 41974 -31442
rect 41174 -31503 41974 -31496
rect 41174 -31600 41974 -31593
rect 41174 -31654 41186 -31600
rect 41962 -31654 41974 -31600
rect 41174 -31661 41974 -31654
rect 41174 -31758 41974 -31751
rect 41174 -31812 41186 -31758
rect 41962 -31812 41974 -31758
rect 41174 -31819 41974 -31812
rect 41174 -31916 41974 -31909
rect 41174 -31970 41186 -31916
rect 41962 -31970 41974 -31916
rect 41174 -31977 41974 -31970
rect 41174 -32074 41974 -32067
rect 41174 -32128 41186 -32074
rect 41962 -32128 41974 -32074
rect 41174 -32135 41974 -32128
rect 41174 -32232 41974 -32225
rect 41174 -32286 41186 -32232
rect 41962 -32286 41974 -32232
rect 41174 -32293 41974 -32286
rect 41174 -32390 41974 -32383
rect 41174 -32444 41186 -32390
rect 41962 -32444 41974 -32390
rect 41174 -32451 41974 -32444
rect 41174 -32548 41974 -32541
rect 41174 -32602 41186 -32548
rect 41962 -32602 41974 -32548
rect 41174 -32609 41974 -32602
rect 41174 -32706 41974 -32699
rect 41174 -32760 41186 -32706
rect 41962 -32760 41974 -32706
rect 41174 -32767 41974 -32760
rect 41174 -32864 41974 -32857
rect 41174 -32918 41186 -32864
rect 41962 -32918 41974 -32864
rect 41174 -32925 41974 -32918
rect 41174 -33022 41974 -33015
rect 41174 -33076 41186 -33022
rect 41962 -33076 41974 -33022
rect 41174 -33083 41974 -33076
rect 41174 -33180 41974 -33173
rect 41174 -33234 41186 -33180
rect 41962 -33234 41974 -33180
rect 41174 -33241 41974 -33234
rect 41174 -33338 41974 -33331
rect 41174 -33392 41186 -33338
rect 41962 -33392 41974 -33338
rect 41174 -33399 41974 -33392
rect 41174 -33496 41974 -33489
rect 41174 -33550 41186 -33496
rect 41962 -33550 41974 -33496
rect 41174 -33557 41974 -33550
rect 41174 -33654 41974 -33647
rect 41174 -33708 41186 -33654
rect 41962 -33708 41974 -33654
rect 41174 -33715 41974 -33708
rect 41174 -33812 41974 -33805
rect 41174 -33866 41186 -33812
rect 41962 -33866 41974 -33812
rect 41174 -33873 41974 -33866
rect 41174 -33970 41974 -33963
rect 41174 -34024 41186 -33970
rect 41962 -34024 41974 -33970
rect 41174 -34031 41974 -34024
rect 41174 -34128 41974 -34121
rect 41174 -34182 41186 -34128
rect 41962 -34182 41974 -34128
rect 41174 -34189 41974 -34182
rect 41174 -34286 41974 -34279
rect 41174 -34340 41186 -34286
rect 41962 -34340 41974 -34286
rect 41174 -34347 41974 -34340
rect 41174 -34444 41974 -34437
rect 41174 -34498 41186 -34444
rect 41962 -34498 41974 -34444
rect 41174 -34505 41974 -34498
rect 41174 -34602 41974 -34595
rect 41174 -34656 41186 -34602
rect 41962 -34656 41974 -34602
rect 41174 -34663 41974 -34656
rect 41174 -34760 41974 -34753
rect 41174 -34814 41186 -34760
rect 41962 -34814 41974 -34760
rect 41174 -34821 41974 -34814
rect 41174 -34918 41974 -34911
rect 41174 -34972 41186 -34918
rect 41962 -34972 41974 -34918
rect 41174 -34979 41974 -34972
rect 41174 -35076 41974 -35069
rect 41174 -35130 41186 -35076
rect 41962 -35130 41974 -35076
rect 41174 -35137 41974 -35130
rect 41174 -35234 41974 -35227
rect 41174 -35288 41186 -35234
rect 41962 -35288 41974 -35234
rect 41174 -35295 41974 -35288
rect 41174 -35392 41974 -35385
rect 41174 -35446 41186 -35392
rect 41962 -35446 41974 -35392
rect 41174 -35453 41974 -35446
rect 41174 -35550 41974 -35543
rect 41174 -35604 41186 -35550
rect 41962 -35604 41974 -35550
rect 41174 -35611 41974 -35604
rect 41174 -35708 41974 -35701
rect 41174 -35762 41186 -35708
rect 41962 -35762 41974 -35708
rect 41174 -35769 41974 -35762
rect 41174 -35866 41974 -35859
rect 41174 -35920 41186 -35866
rect 41962 -35920 41974 -35866
rect 41174 -35927 41974 -35920
rect 41174 -36024 41974 -36017
rect 41174 -36078 41186 -36024
rect 41962 -36078 41974 -36024
rect 41174 -36085 41974 -36078
rect 41174 -36182 41974 -36175
rect 41174 -36236 41186 -36182
rect 41962 -36236 41974 -36182
rect 41174 -36243 41974 -36236
rect 41174 -36340 41974 -36333
rect 41174 -36394 41186 -36340
rect 41962 -36394 41974 -36340
rect 41174 -36401 41974 -36394
rect 41174 -36498 41974 -36491
rect 41174 -36552 41186 -36498
rect 41962 -36552 41974 -36498
rect 41174 -36559 41974 -36552
rect 41174 -36656 41974 -36649
rect 41174 -36710 41186 -36656
rect 41962 -36710 41974 -36656
rect 41174 -36717 41974 -36710
rect 41174 -36814 41974 -36807
rect 41174 -36868 41186 -36814
rect 41962 -36868 41974 -36814
rect 41174 -36875 41974 -36868
rect 41174 -36972 41974 -36965
rect 41174 -37026 41186 -36972
rect 41962 -37026 41974 -36972
rect 41174 -37033 41974 -37026
rect 41174 -37130 41974 -37123
rect 41174 -37184 41186 -37130
rect 41962 -37184 41974 -37130
rect 41174 -37191 41974 -37184
rect 41174 -37288 41974 -37281
rect 41174 -37342 41186 -37288
rect 41962 -37342 41974 -37288
rect 41174 -37349 41974 -37342
rect 41174 -37446 41974 -37439
rect 41174 -37500 41186 -37446
rect 41962 -37500 41974 -37446
rect 41174 -37507 41974 -37500
rect 41174 -37604 41974 -37597
rect 41174 -37658 41186 -37604
rect 41962 -37658 41974 -37604
rect 41174 -37665 41974 -37658
rect 41174 -37762 41974 -37755
rect 41174 -37816 41186 -37762
rect 41962 -37816 41974 -37762
rect 41174 -37823 41974 -37816
rect 41174 -37920 41974 -37913
rect 41174 -37974 41186 -37920
rect 41962 -37974 41974 -37920
rect 41174 -37981 41974 -37974
rect 41174 -38078 41974 -38071
rect 41174 -38132 41186 -38078
rect 41962 -38132 41974 -38078
rect 41174 -38139 41974 -38132
rect 41174 -38236 41974 -38229
rect 41174 -38290 41186 -38236
rect 41962 -38290 41974 -38236
rect 41174 -38297 41974 -38290
rect 41174 -38394 41974 -38387
rect 41174 -38448 41186 -38394
rect 41962 -38448 41974 -38394
rect 41174 -38455 41974 -38448
rect 41174 -38552 41974 -38545
rect 42006 -38550 42062 -26023
rect 41174 -38606 41186 -38552
rect 41962 -38606 41974 -38552
rect 41174 -38613 41974 -38606
rect 42138 -38684 42196 -25834
rect 40952 -38742 42196 -38684
rect 3771 -44081 11640 -43796
rect 368 -45580 3619 -45524
rect 368 -45771 424 -45580
rect 606 -45656 2112 -45649
rect 606 -45685 642 -45656
rect 1967 -45685 2112 -45656
rect 606 -45719 630 -45685
rect 1980 -45719 2112 -45685
rect 606 -45729 642 -45719
rect 1967 -45729 2112 -45719
rect 606 -45735 2112 -45729
rect 368 -45827 822 -45771
rect 2022 -45781 2112 -45735
rect 368 -46898 424 -45827
rect 2022 -45868 2042 -45781
rect 498 -45874 694 -45868
rect 360 -46912 432 -46898
rect 360 -46968 368 -46912
rect 424 -46968 432 -46912
rect 360 -46974 432 -46968
rect 498 -46955 534 -45874
rect 568 -45875 694 -45874
rect 568 -46862 639 -45875
rect 692 -46862 694 -45875
rect 568 -46868 694 -46862
rect 764 -45875 822 -45868
rect 764 -46862 767 -45875
rect 820 -46862 822 -45875
rect 764 -46868 822 -46862
rect 892 -45875 950 -45868
rect 892 -46862 895 -45875
rect 948 -46862 950 -45875
rect 892 -46868 950 -46862
rect 1020 -45875 1078 -45868
rect 1020 -46862 1023 -45875
rect 1076 -46862 1078 -45875
rect 1020 -46868 1078 -46862
rect 1148 -45875 1206 -45868
rect 1148 -46862 1151 -45875
rect 1204 -46862 1206 -45875
rect 1148 -46868 1206 -46862
rect 1276 -45875 1334 -45868
rect 1276 -46862 1279 -45875
rect 1332 -46862 1334 -45875
rect 1276 -46868 1334 -46862
rect 1404 -45875 1462 -45868
rect 1404 -46862 1407 -45875
rect 1460 -46862 1462 -45875
rect 1404 -46868 1462 -46862
rect 1532 -45875 1590 -45868
rect 1532 -46862 1535 -45875
rect 1588 -46862 1590 -45875
rect 1532 -46868 1590 -46862
rect 1660 -45875 1718 -45868
rect 1660 -46862 1663 -45875
rect 1716 -46862 1718 -45875
rect 1660 -46868 1718 -46862
rect 1788 -45875 1846 -45868
rect 1788 -46862 1791 -45875
rect 1844 -46862 1846 -45875
rect 1788 -46868 1846 -46862
rect 1916 -45875 2042 -45868
rect 1916 -46862 1919 -45875
rect 1972 -46862 2042 -45875
rect 1916 -46868 2042 -46862
rect 568 -46955 578 -46868
rect 498 -47008 578 -46955
rect 614 -46909 682 -46903
rect 1904 -46907 1989 -46901
rect 1904 -46909 1911 -46907
rect 614 -46965 620 -46909
rect 676 -46965 946 -46909
rect 1896 -46960 1911 -46909
rect 1983 -46960 1989 -46907
rect 1896 -46965 1989 -46960
rect 2022 -46955 2042 -46868
rect 2076 -46955 2112 -45781
rect 614 -46971 682 -46965
rect 2022 -47008 2112 -46955
rect 498 -47017 2112 -47008
rect 498 -47051 630 -47017
rect 1980 -47051 2112 -47017
rect 498 -47087 2112 -47051
rect 498 -47341 602 -47087
rect 2008 -47341 2112 -47087
rect 498 -47377 2112 -47341
rect 498 -47411 630 -47377
rect 1980 -47411 2112 -47377
rect 498 -47427 2112 -47411
rect 498 -47473 588 -47427
rect 498 -48647 534 -47473
rect 568 -48647 588 -47473
rect 1902 -47461 1987 -47455
rect 1902 -47514 1909 -47461
rect 1981 -47514 1987 -47461
rect 1902 -47519 1987 -47514
rect 2022 -47473 2112 -47427
rect 636 -47567 694 -47560
rect 636 -48554 639 -47567
rect 692 -48554 694 -47567
rect 636 -48560 694 -48554
rect 764 -47567 822 -47560
rect 764 -48554 767 -47567
rect 820 -48554 822 -47567
rect 764 -48560 822 -48554
rect 892 -47567 950 -47560
rect 892 -48554 895 -47567
rect 948 -48554 950 -47567
rect 892 -48560 950 -48554
rect 1020 -47567 1078 -47560
rect 1020 -48554 1023 -47567
rect 1076 -48554 1078 -47567
rect 1020 -48560 1078 -48554
rect 1148 -47567 1206 -47560
rect 1148 -48554 1151 -47567
rect 1204 -48554 1206 -47567
rect 1148 -48560 1206 -48554
rect 1276 -47567 1334 -47560
rect 1276 -48554 1279 -47567
rect 1332 -48554 1334 -47567
rect 1276 -48560 1334 -48554
rect 1404 -47567 1462 -47560
rect 1404 -48554 1407 -47567
rect 1460 -48554 1462 -47567
rect 1404 -48560 1462 -48554
rect 1532 -47567 1590 -47560
rect 1532 -48554 1535 -47567
rect 1588 -48554 1590 -47567
rect 1532 -48560 1590 -48554
rect 1660 -47567 1718 -47560
rect 1660 -48554 1663 -47567
rect 1716 -48554 1718 -47567
rect 1660 -48560 1718 -48554
rect 1788 -47567 1846 -47560
rect 1788 -48554 1791 -47567
rect 1844 -48554 1846 -47567
rect 1788 -48560 1846 -48554
rect 1916 -47567 1974 -47560
rect 1916 -48554 1919 -47567
rect 1972 -48554 1974 -47567
rect 1916 -48560 1974 -48554
rect 498 -48693 588 -48647
rect 498 -48709 1227 -48693
rect 498 -48743 630 -48709
rect 1221 -48743 1227 -48709
rect 498 -48779 1227 -48743
rect 1269 -48822 1339 -48629
rect 2022 -48647 2042 -47473
rect 2076 -48647 2112 -47473
rect 2022 -48693 2112 -48647
rect 1367 -48709 2112 -48693
rect 1367 -48743 1373 -48709
rect 1980 -48743 2112 -48709
rect 1367 -48779 2112 -48743
rect 2214 -46340 2802 -46263
rect 2214 -46395 2304 -46340
rect 2834 -46385 2890 -45580
rect 3563 -45863 3619 -45580
rect 3541 -45888 3646 -45863
rect 3541 -45944 3563 -45888
rect 3619 -45944 3646 -45888
rect 3541 -45961 3646 -45944
rect 2919 -46340 3508 -46263
rect 2214 -46951 2250 -46395
rect 2284 -46951 2304 -46395
rect 2492 -46441 3326 -46385
rect 3432 -46395 3508 -46340
rect 2348 -46867 2354 -46473
rect 2408 -46867 2414 -46473
rect 2348 -46873 2414 -46867
rect 2444 -46867 2450 -46473
rect 2504 -46867 2510 -46473
rect 2444 -46873 2510 -46867
rect 2540 -46867 2546 -46473
rect 2600 -46867 2606 -46473
rect 2540 -46873 2606 -46867
rect 2636 -46867 2642 -46473
rect 2696 -46867 2702 -46473
rect 2636 -46873 2702 -46867
rect 2732 -46867 2738 -46473
rect 2792 -46867 2798 -46473
rect 2732 -46873 2798 -46867
rect 2828 -46867 2834 -46473
rect 2888 -46867 2894 -46473
rect 2828 -46873 2894 -46867
rect 2924 -46867 2930 -46473
rect 2984 -46867 2990 -46473
rect 2924 -46873 2990 -46867
rect 3020 -46867 3026 -46473
rect 3080 -46867 3086 -46473
rect 3020 -46873 3086 -46867
rect 3116 -46867 3122 -46473
rect 3176 -46867 3182 -46473
rect 3116 -46873 3182 -46867
rect 3212 -46867 3218 -46473
rect 3272 -46867 3278 -46473
rect 3212 -46873 3278 -46867
rect 3308 -46867 3314 -46473
rect 3368 -46867 3374 -46473
rect 3308 -46873 3374 -46867
rect 2214 -47007 2304 -46951
rect 2332 -46905 2396 -46901
rect 3314 -46905 3396 -46901
rect 2332 -46907 3396 -46905
rect 2332 -46908 3320 -46907
rect 2332 -46961 2338 -46908
rect 2390 -46961 3320 -46908
rect 2332 -46963 3320 -46961
rect 3390 -46963 3396 -46907
rect 2332 -46966 3396 -46963
rect 2332 -46967 2396 -46966
rect 3314 -46971 3396 -46966
rect 3432 -46951 3438 -46395
rect 3472 -46951 3508 -46395
rect 3432 -47007 3508 -46951
rect 2214 -47013 3508 -47007
rect 2214 -47047 2346 -47013
rect 3376 -47047 3508 -47013
rect 2214 -47083 3508 -47047
rect 2214 -47341 2356 -47083
rect 3366 -47341 3508 -47083
rect 2214 -47426 3508 -47341
rect 2214 -47551 2296 -47426
rect 2324 -47460 2409 -47454
rect 2324 -47513 2331 -47460
rect 2403 -47463 2409 -47460
rect 2403 -47513 2787 -47463
rect 2324 -47519 2787 -47513
rect 2214 -48141 2304 -47551
rect 2731 -47821 2787 -47519
rect 3312 -47776 3387 -47757
rect 3312 -47821 3322 -47776
rect 2731 -47877 3322 -47821
rect 2214 -48177 2657 -48141
rect 2214 -48211 2346 -48177
rect 2621 -48211 2657 -48177
rect 2214 -48229 2657 -48211
rect 2214 -48273 2304 -48229
rect 2731 -48263 2787 -47877
rect 3312 -47909 3322 -47877
rect 3374 -47909 3387 -47776
rect 3312 -47923 3387 -47909
rect 3418 -48141 3508 -47426
rect 3771 -47726 4056 -44081
rect 3079 -48177 3508 -48141
rect 3079 -48211 3101 -48177
rect 3376 -48211 3508 -48177
rect 3079 -48229 3508 -48211
rect 2214 -48629 2250 -48273
rect 2284 -48351 2304 -48273
rect 2492 -48319 3326 -48263
rect 3418 -48273 3508 -48229
rect 3418 -48351 3438 -48273
rect 2284 -48545 2354 -48351
rect 2408 -48545 2414 -48351
rect 2284 -48551 2414 -48545
rect 2444 -48545 2450 -48351
rect 2504 -48545 2510 -48351
rect 2444 -48551 2510 -48545
rect 2540 -48545 2546 -48351
rect 2600 -48545 2606 -48351
rect 2540 -48551 2606 -48545
rect 2636 -48545 2642 -48351
rect 2696 -48545 2702 -48351
rect 2636 -48551 2702 -48545
rect 2732 -48545 2738 -48351
rect 2792 -48545 2798 -48351
rect 2732 -48551 2798 -48545
rect 2828 -48545 2834 -48351
rect 2888 -48545 2894 -48351
rect 2828 -48551 2894 -48545
rect 2924 -48545 2930 -48351
rect 2984 -48545 2990 -48351
rect 2924 -48551 2990 -48545
rect 3020 -48545 3026 -48351
rect 3080 -48545 3086 -48351
rect 3020 -48551 3086 -48545
rect 3116 -48545 3122 -48351
rect 3176 -48545 3182 -48351
rect 3116 -48551 3182 -48545
rect 3212 -48545 3218 -48351
rect 3272 -48545 3278 -48351
rect 3212 -48551 3278 -48545
rect 3308 -48545 3314 -48351
rect 3368 -48545 3438 -48351
rect 3308 -48551 3438 -48545
rect 2284 -48629 2304 -48551
rect 2214 -48671 2304 -48629
rect 2396 -48639 3230 -48583
rect 3418 -48629 3438 -48551
rect 3472 -48629 3508 -48273
rect 2214 -48677 2798 -48671
rect 2214 -48691 2354 -48677
rect 2214 -48725 2346 -48691
rect 2214 -48755 2354 -48725
rect 2792 -48755 2798 -48677
rect 2214 -48761 2798 -48755
rect 2826 -48822 2896 -48639
rect 3418 -48671 3508 -48629
rect 2924 -48677 3508 -48671
rect 2924 -48755 2930 -48677
rect 3368 -48691 3508 -48677
rect 3376 -48725 3508 -48691
rect 3368 -48755 3508 -48725
rect 2924 -48761 3508 -48755
rect 3567 -47770 4056 -47726
rect 3567 -47909 3683 -47770
rect 3822 -47909 4056 -47770
rect 3567 -48047 4056 -47909
rect 3567 -48822 3637 -48047
rect -6172 -49150 -5411 -48864
rect 1269 -48892 3637 -48822
rect 2348 -48988 3374 -48963
rect 2348 -49150 2391 -48988
rect 3339 -49150 3374 -48988
rect -6172 -49536 -6013 -49150
rect -5627 -49536 3374 -49150
rect -6172 -49739 -5411 -49536
rect -1558 -51813 -1172 -49536
rect 41551 -51813 41937 -38742
rect -1558 -52199 41937 -51813
<< via1 >>
rect 12686 739 12778 831
rect -196 540 -98 638
rect 211 233 297 239
rect 211 159 219 233
rect 219 159 294 233
rect 294 159 297 233
rect 211 153 297 159
rect 377 233 467 246
rect 377 167 401 233
rect 401 167 467 233
rect 377 160 467 167
rect 517 233 607 259
rect 517 165 581 233
rect 581 165 607 233
rect 885 267 937 346
rect 885 165 892 267
rect 892 165 926 267
rect 926 165 937 267
rect 885 162 937 165
rect 1062 251 1137 257
rect 1062 185 1068 251
rect 1068 185 1133 251
rect 1133 185 1137 251
rect 1062 179 1137 185
rect 3298 177 3392 279
rect 3573 313 3589 346
rect 3589 313 3623 346
rect 3623 313 3625 346
rect 3573 267 3625 313
rect 3573 165 3580 267
rect 3580 165 3614 267
rect 3614 165 3625 267
rect 3573 162 3625 165
rect 3750 251 3825 257
rect 3750 185 3756 251
rect 3756 185 3821 251
rect 3821 185 3825 251
rect 3750 179 3825 185
rect 5986 177 6080 279
rect 6261 313 6277 346
rect 6277 313 6311 346
rect 6311 313 6313 346
rect 6261 267 6313 313
rect 6261 165 6268 267
rect 6268 165 6302 267
rect 6302 165 6313 267
rect 6261 162 6313 165
rect 6438 251 6513 257
rect 6438 185 6444 251
rect 6444 185 6509 251
rect 6509 185 6513 251
rect 6438 179 6513 185
rect 8674 177 8768 279
rect 8949 313 8965 346
rect 8965 313 8999 346
rect 8999 313 9001 346
rect 8949 267 9001 313
rect 8949 165 8956 267
rect 8956 165 8990 267
rect 8990 165 9001 267
rect 8949 162 9001 165
rect 9126 251 9201 257
rect 9126 185 9132 251
rect 9132 185 9197 251
rect 9197 185 9201 251
rect 9126 179 9201 185
rect 11362 177 11456 279
rect -5966 -552 -5627 -213
rect -196 -792 -98 -694
rect 2615 -1012 2865 -893
rect 5303 -1002 5553 -893
rect 8001 -1007 8222 -903
rect 10686 -1006 10902 -903
rect 3298 -1189 3565 -1058
rect 5986 -1189 6253 -1073
rect 8692 -1159 8926 -1072
rect 11378 -1166 11608 -1078
rect 19140 400 19460 720
rect 19171 -206 19429 52
rect 19302 -802 19354 -615
rect 19206 -933 19286 -862
rect 12873 -1219 12943 -1149
rect 18779 -1648 18944 -1483
rect 19217 -1414 19298 -1347
rect 19315 -1650 19367 -1466
rect -196 -2124 -98 -2026
rect 14187 -2133 14277 -2043
rect 2599 -2710 2883 -2426
rect 5287 -2710 5571 -2426
rect 7975 -2710 8259 -2426
rect 10663 -2710 10947 -2426
rect 12320 -2630 12736 -2572
rect 3292 -3290 3576 -3006
rect 642 -3685 1967 -3656
rect 642 -3719 1967 -3685
rect 642 -3729 1967 -3719
rect 368 -4968 424 -4912
rect 639 -4862 692 -3875
rect 767 -4862 820 -3875
rect 895 -4862 948 -3875
rect 1023 -4862 1076 -3875
rect 1151 -4862 1204 -3875
rect 1279 -4862 1332 -3875
rect 1407 -4862 1460 -3875
rect 1535 -4862 1588 -3875
rect 1663 -4862 1716 -3875
rect 1791 -4862 1844 -3875
rect 1919 -4862 1972 -3875
rect 620 -4965 676 -4909
rect 1911 -4960 1983 -4907
rect 1909 -5514 1981 -5461
rect 639 -6554 692 -5567
rect 767 -6554 820 -5567
rect 895 -6554 948 -5567
rect 1023 -6554 1076 -5567
rect 1151 -6554 1204 -5567
rect 1279 -6554 1332 -5567
rect 1407 -6554 1460 -5567
rect 1535 -6554 1588 -5567
rect 1663 -6554 1716 -5567
rect 1791 -6554 1844 -5567
rect 1919 -6554 1972 -5567
rect 3563 -3944 3619 -3888
rect 2354 -4867 2408 -4473
rect 2450 -4867 2504 -4473
rect 2546 -4867 2600 -4473
rect 2642 -4867 2696 -4473
rect 2738 -4867 2792 -4473
rect 2834 -4867 2888 -4473
rect 2930 -4867 2984 -4473
rect 3026 -4867 3080 -4473
rect 3122 -4867 3176 -4473
rect 3218 -4867 3272 -4473
rect 3314 -4867 3368 -4473
rect 2338 -4961 2390 -4908
rect 3320 -4963 3390 -4907
rect 2331 -5513 2403 -5460
rect 3322 -5909 3374 -5776
rect 2354 -6545 2408 -6351
rect 2450 -6545 2504 -6351
rect 2546 -6545 2600 -6351
rect 2642 -6545 2696 -6351
rect 2738 -6545 2792 -6351
rect 2834 -6545 2888 -6351
rect 2930 -6545 2984 -6351
rect 3026 -6545 3080 -6351
rect 3122 -6545 3176 -6351
rect 3218 -6545 3272 -6351
rect 3314 -6545 3368 -6351
rect 2354 -6691 2792 -6677
rect 2354 -6725 2792 -6691
rect 2354 -6755 2792 -6725
rect 2930 -6691 3368 -6677
rect 2930 -6725 3368 -6691
rect 2930 -6755 3368 -6725
rect 3683 -5909 3822 -5770
rect 2391 -7150 3339 -6988
rect -6013 -7536 -5627 -7150
rect 5980 -3009 6264 -2725
rect 642 -17685 1967 -17656
rect 642 -17719 1967 -17685
rect 642 -17729 1967 -17719
rect 368 -18968 424 -18912
rect 639 -18862 692 -17875
rect 767 -18862 820 -17875
rect 895 -18862 948 -17875
rect 1023 -18862 1076 -17875
rect 1151 -18862 1204 -17875
rect 1279 -18862 1332 -17875
rect 1407 -18862 1460 -17875
rect 1535 -18862 1588 -17875
rect 1663 -18862 1716 -17875
rect 1791 -18862 1844 -17875
rect 1919 -18862 1972 -17875
rect 620 -18965 676 -18909
rect 1911 -18960 1983 -18907
rect 1909 -19514 1981 -19461
rect 639 -20554 692 -19567
rect 767 -20554 820 -19567
rect 895 -20554 948 -19567
rect 1023 -20554 1076 -19567
rect 1151 -20554 1204 -19567
rect 1279 -20554 1332 -19567
rect 1407 -20554 1460 -19567
rect 1535 -20554 1588 -19567
rect 1663 -20554 1716 -19567
rect 1791 -20554 1844 -19567
rect 1919 -20554 1972 -19567
rect 3563 -17944 3619 -17888
rect 2354 -18867 2408 -18473
rect 2450 -18867 2504 -18473
rect 2546 -18867 2600 -18473
rect 2642 -18867 2696 -18473
rect 2738 -18867 2792 -18473
rect 2834 -18867 2888 -18473
rect 2930 -18867 2984 -18473
rect 3026 -18867 3080 -18473
rect 3122 -18867 3176 -18473
rect 3218 -18867 3272 -18473
rect 3314 -18867 3368 -18473
rect 2338 -18961 2390 -18908
rect 3320 -18963 3390 -18907
rect 2331 -19513 2403 -19460
rect 3322 -19909 3374 -19776
rect 2354 -20545 2408 -20351
rect 2450 -20545 2504 -20351
rect 2546 -20545 2600 -20351
rect 2642 -20545 2696 -20351
rect 2738 -20545 2792 -20351
rect 2834 -20545 2888 -20351
rect 2930 -20545 2984 -20351
rect 3026 -20545 3080 -20351
rect 3122 -20545 3176 -20351
rect 3218 -20545 3272 -20351
rect 3314 -20545 3368 -20351
rect 2354 -20691 2792 -20677
rect 2354 -20725 2792 -20691
rect 2354 -20755 2792 -20725
rect 2930 -20691 3368 -20677
rect 2930 -20725 3368 -20691
rect 2930 -20755 3368 -20725
rect 3683 -19909 3822 -19770
rect 2391 -21150 3339 -20988
rect -6013 -21536 -5627 -21150
rect 8668 -3316 8952 -3032
rect 642 -31685 1967 -31656
rect 642 -31719 1967 -31685
rect 642 -31729 1967 -31719
rect 368 -32968 424 -32912
rect 639 -32862 692 -31875
rect 767 -32862 820 -31875
rect 895 -32862 948 -31875
rect 1023 -32862 1076 -31875
rect 1151 -32862 1204 -31875
rect 1279 -32862 1332 -31875
rect 1407 -32862 1460 -31875
rect 1535 -32862 1588 -31875
rect 1663 -32862 1716 -31875
rect 1791 -32862 1844 -31875
rect 1919 -32862 1972 -31875
rect 620 -32965 676 -32909
rect 1911 -32960 1983 -32907
rect 1909 -33514 1981 -33461
rect 639 -34554 692 -33567
rect 767 -34554 820 -33567
rect 895 -34554 948 -33567
rect 1023 -34554 1076 -33567
rect 1151 -34554 1204 -33567
rect 1279 -34554 1332 -33567
rect 1407 -34554 1460 -33567
rect 1535 -34554 1588 -33567
rect 1663 -34554 1716 -33567
rect 1791 -34554 1844 -33567
rect 1919 -34554 1972 -33567
rect 3563 -31944 3619 -31888
rect 2354 -32867 2408 -32473
rect 2450 -32867 2504 -32473
rect 2546 -32867 2600 -32473
rect 2642 -32867 2696 -32473
rect 2738 -32867 2792 -32473
rect 2834 -32867 2888 -32473
rect 2930 -32867 2984 -32473
rect 3026 -32867 3080 -32473
rect 3122 -32867 3176 -32473
rect 3218 -32867 3272 -32473
rect 3314 -32867 3368 -32473
rect 2338 -32961 2390 -32908
rect 3320 -32963 3390 -32907
rect 2331 -33513 2403 -33460
rect 3322 -33909 3374 -33776
rect 2354 -34545 2408 -34351
rect 2450 -34545 2504 -34351
rect 2546 -34545 2600 -34351
rect 2642 -34545 2696 -34351
rect 2738 -34545 2792 -34351
rect 2834 -34545 2888 -34351
rect 2930 -34545 2984 -34351
rect 3026 -34545 3080 -34351
rect 3122 -34545 3176 -34351
rect 3218 -34545 3272 -34351
rect 3314 -34545 3368 -34351
rect 2354 -34691 2792 -34677
rect 2354 -34725 2792 -34691
rect 2354 -34755 2792 -34725
rect 2930 -34691 3368 -34677
rect 2930 -34725 3368 -34691
rect 2930 -34755 3368 -34725
rect 3683 -33909 3822 -33770
rect 2391 -35150 3339 -34988
rect -6013 -35536 -5627 -35150
rect 13088 -2630 13504 -2572
rect 13850 -2630 14266 -2572
rect 11356 -3476 11640 -3192
rect 41203 -11921 41979 -11867
rect 42050 -11916 42114 -11849
rect 41203 -12079 41979 -12025
rect 41203 -12237 41979 -12183
rect 41203 -12395 41979 -12341
rect 41203 -12553 41979 -12499
rect 41203 -12711 41979 -12657
rect 41203 -12869 41979 -12815
rect 41203 -13027 41979 -12973
rect 41203 -13185 41979 -13131
rect 41203 -13343 41979 -13289
rect 41203 -13501 41979 -13447
rect 41203 -13659 41979 -13605
rect 41203 -13817 41979 -13763
rect 41203 -13975 41979 -13921
rect 41203 -14133 41979 -14079
rect 41203 -14291 41979 -14237
rect 41203 -14449 41979 -14395
rect 41203 -14607 41979 -14553
rect 41203 -14765 41979 -14711
rect 41203 -14923 41979 -14869
rect 41203 -15081 41979 -15027
rect 41203 -15239 41979 -15185
rect 41203 -15397 41979 -15343
rect 41203 -15555 41979 -15501
rect 41203 -15713 41979 -15659
rect 41203 -15871 41979 -15817
rect 41203 -16029 41979 -15975
rect 41203 -16187 41979 -16133
rect 41203 -16345 41979 -16291
rect 41203 -16503 41979 -16449
rect 41203 -16661 41979 -16607
rect 41203 -16819 41979 -16765
rect 41203 -16977 41979 -16923
rect 41203 -17135 41979 -17081
rect 41203 -17293 41979 -17239
rect 41203 -17451 41979 -17397
rect 41203 -17609 41979 -17555
rect 41203 -17767 41979 -17713
rect 41203 -17925 41979 -17871
rect 41203 -18083 41979 -18029
rect 41203 -18241 41979 -18187
rect 41203 -18399 41979 -18345
rect 41203 -18557 41979 -18503
rect 41203 -18715 41979 -18661
rect 41203 -18873 41979 -18819
rect 41203 -19031 41979 -18977
rect 41203 -19189 41979 -19135
rect 41203 -19347 41979 -19293
rect 41203 -19505 41979 -19451
rect 41203 -19663 41979 -19609
rect 41203 -19821 41979 -19767
rect 41203 -19979 41979 -19925
rect 41203 -20137 41979 -20083
rect 41203 -20295 41979 -20241
rect 41203 -20453 41979 -20399
rect 41203 -20611 41979 -20557
rect 41203 -20769 41979 -20715
rect 41203 -20927 41979 -20873
rect 41203 -21085 41979 -21031
rect 41203 -21243 41979 -21189
rect 41203 -21401 41979 -21347
rect 41203 -21559 41979 -21505
rect 41203 -21717 41979 -21663
rect 41203 -21875 41979 -21821
rect 41203 -22033 41979 -21979
rect 41203 -22191 41979 -22137
rect 41203 -22349 41979 -22295
rect 41203 -22507 41979 -22453
rect 41203 -22665 41979 -22611
rect 41203 -22823 41979 -22769
rect 41203 -22981 41979 -22927
rect 41203 -23139 41979 -23085
rect 41203 -23297 41979 -23243
rect 41203 -23455 41979 -23401
rect 41203 -23613 41979 -23559
rect 41203 -23771 41979 -23717
rect 41203 -23929 41979 -23875
rect 41203 -24087 41979 -24033
rect 41203 -24245 41979 -24191
rect 41203 -24403 41979 -24349
rect 41203 -24561 41979 -24507
rect 41186 -25966 41962 -25912
rect 41053 -26151 41128 -26056
rect 42014 -26014 42098 -25946
rect 41186 -26124 41962 -26070
rect 41186 -26282 41962 -26228
rect 41186 -26440 41962 -26386
rect 41186 -26598 41962 -26544
rect 41186 -26756 41962 -26702
rect 41186 -26914 41962 -26860
rect 41186 -27072 41962 -27018
rect 41186 -27230 41962 -27176
rect 41186 -27388 41962 -27334
rect 41186 -27546 41962 -27492
rect 41186 -27704 41962 -27650
rect 41186 -27862 41962 -27808
rect 41186 -28020 41962 -27966
rect 41186 -28178 41962 -28124
rect 41186 -28336 41962 -28282
rect 41186 -28494 41962 -28440
rect 41186 -28652 41962 -28598
rect 41186 -28810 41962 -28756
rect 41186 -28968 41962 -28914
rect 41186 -29126 41962 -29072
rect 41186 -29284 41962 -29230
rect 41186 -29442 41962 -29388
rect 41186 -29600 41962 -29546
rect 41186 -29758 41962 -29704
rect 41186 -29916 41962 -29862
rect 41186 -30074 41962 -30020
rect 41186 -30232 41962 -30178
rect 41186 -30390 41962 -30336
rect 41186 -30548 41962 -30494
rect 41186 -30706 41962 -30652
rect 41186 -30864 41962 -30810
rect 41186 -31022 41962 -30968
rect 41186 -31180 41962 -31126
rect 41186 -31338 41962 -31284
rect 41186 -31496 41962 -31442
rect 41186 -31654 41962 -31600
rect 41186 -31812 41962 -31758
rect 41186 -31970 41962 -31916
rect 41186 -32128 41962 -32074
rect 41186 -32286 41962 -32232
rect 41186 -32444 41962 -32390
rect 41186 -32602 41962 -32548
rect 41186 -32760 41962 -32706
rect 41186 -32918 41962 -32864
rect 41186 -33076 41962 -33022
rect 41186 -33234 41962 -33180
rect 41186 -33392 41962 -33338
rect 41186 -33550 41962 -33496
rect 41186 -33708 41962 -33654
rect 41186 -33866 41962 -33812
rect 41186 -34024 41962 -33970
rect 41186 -34182 41962 -34128
rect 41186 -34340 41962 -34286
rect 41186 -34498 41962 -34444
rect 41186 -34656 41962 -34602
rect 41186 -34814 41962 -34760
rect 41186 -34972 41962 -34918
rect 41186 -35130 41962 -35076
rect 41186 -35288 41962 -35234
rect 41186 -35446 41962 -35392
rect 41186 -35604 41962 -35550
rect 41186 -35762 41962 -35708
rect 41186 -35920 41962 -35866
rect 41186 -36078 41962 -36024
rect 41186 -36236 41962 -36182
rect 41186 -36394 41962 -36340
rect 41186 -36552 41962 -36498
rect 41186 -36710 41962 -36656
rect 41186 -36868 41962 -36814
rect 41186 -37026 41962 -36972
rect 41186 -37184 41962 -37130
rect 41186 -37342 41962 -37288
rect 41186 -37500 41962 -37446
rect 41186 -37658 41962 -37604
rect 41186 -37816 41962 -37762
rect 41186 -37974 41962 -37920
rect 41186 -38132 41962 -38078
rect 41186 -38290 41962 -38236
rect 41186 -38448 41962 -38394
rect 41186 -38606 41962 -38552
rect 642 -45685 1967 -45656
rect 642 -45719 1967 -45685
rect 642 -45729 1967 -45719
rect 368 -46968 424 -46912
rect 639 -46862 692 -45875
rect 767 -46862 820 -45875
rect 895 -46862 948 -45875
rect 1023 -46862 1076 -45875
rect 1151 -46862 1204 -45875
rect 1279 -46862 1332 -45875
rect 1407 -46862 1460 -45875
rect 1535 -46862 1588 -45875
rect 1663 -46862 1716 -45875
rect 1791 -46862 1844 -45875
rect 1919 -46862 1972 -45875
rect 620 -46965 676 -46909
rect 1911 -46960 1983 -46907
rect 1909 -47514 1981 -47461
rect 639 -48554 692 -47567
rect 767 -48554 820 -47567
rect 895 -48554 948 -47567
rect 1023 -48554 1076 -47567
rect 1151 -48554 1204 -47567
rect 1279 -48554 1332 -47567
rect 1407 -48554 1460 -47567
rect 1535 -48554 1588 -47567
rect 1663 -48554 1716 -47567
rect 1791 -48554 1844 -47567
rect 1919 -48554 1972 -47567
rect 3563 -45944 3619 -45888
rect 2354 -46867 2408 -46473
rect 2450 -46867 2504 -46473
rect 2546 -46867 2600 -46473
rect 2642 -46867 2696 -46473
rect 2738 -46867 2792 -46473
rect 2834 -46867 2888 -46473
rect 2930 -46867 2984 -46473
rect 3026 -46867 3080 -46473
rect 3122 -46867 3176 -46473
rect 3218 -46867 3272 -46473
rect 3314 -46867 3368 -46473
rect 2338 -46961 2390 -46908
rect 3320 -46963 3390 -46907
rect 2331 -47513 2403 -47460
rect 3322 -47909 3374 -47776
rect 2354 -48545 2408 -48351
rect 2450 -48545 2504 -48351
rect 2546 -48545 2600 -48351
rect 2642 -48545 2696 -48351
rect 2738 -48545 2792 -48351
rect 2834 -48545 2888 -48351
rect 2930 -48545 2984 -48351
rect 3026 -48545 3080 -48351
rect 3122 -48545 3176 -48351
rect 3218 -48545 3272 -48351
rect 3314 -48545 3368 -48351
rect 2354 -48691 2792 -48677
rect 2354 -48725 2792 -48691
rect 2354 -48755 2792 -48725
rect 2930 -48691 3368 -48677
rect 2930 -48725 3368 -48691
rect 2930 -48755 3368 -48725
rect 3683 -47909 3822 -47770
rect 2391 -49150 3339 -48988
rect -6013 -49536 -5627 -49150
<< metal2 >>
rect -4072 2059 -3400 2092
rect -4072 1487 -4014 2059
rect -3442 1487 17110 2059
rect -4072 1429 -3400 1487
rect 205 969 8773 1067
rect -253 638 -32 655
rect -253 540 -196 638
rect -98 540 -32 638
rect -6127 -213 -5411 -70
rect -6127 -552 -5966 -213
rect -5627 -552 -5411 -213
rect -6127 -683 -5411 -552
rect -253 -694 -32 540
rect 205 239 303 969
rect 205 153 211 239
rect 297 153 303 239
rect 371 823 6085 925
rect 371 246 473 823
rect 371 160 377 246
rect 467 160 473 246
rect 371 154 473 160
rect 509 681 3397 786
rect 509 259 614 681
rect 509 165 517 259
rect 607 165 614 259
rect 509 158 614 165
rect 879 346 947 353
rect 879 162 885 346
rect 937 162 947 346
rect 3292 291 3397 681
rect 3567 346 3635 353
rect 3292 279 3398 291
rect 205 147 303 153
rect 879 -295 947 162
rect 1056 257 1145 263
rect 1056 179 1062 257
rect 1137 179 1145 257
rect 1056 -146 1145 179
rect 1056 -217 1065 -146
rect 1136 -217 1145 -146
rect 1056 -226 1145 -217
rect 3292 177 3298 279
rect 3392 177 3398 279
rect 868 -306 958 -295
rect 868 -374 879 -306
rect 947 -374 958 -306
rect 868 -385 958 -374
rect -253 -792 -196 -694
rect -98 -792 -32 -694
rect -253 -2026 -32 -792
rect -253 -2124 -196 -2026
rect -98 -2124 -32 -2026
rect -4155 -2876 -3272 -2759
rect -253 -2876 -32 -2124
rect 2599 -893 2883 -879
rect 2599 -1012 2615 -893
rect 2865 -1012 2883 -893
rect 2599 -2426 2883 -1012
rect 2599 -2716 2883 -2710
rect 3292 -1053 3398 177
rect 3567 162 3573 346
rect 3625 162 3635 346
rect 5980 291 6085 823
rect 6255 346 6323 353
rect 5980 279 6086 291
rect 3567 -295 3635 162
rect 3744 257 3833 263
rect 3744 179 3750 257
rect 3825 179 3833 257
rect 3744 -146 3833 179
rect 5981 177 5986 279
rect 6080 177 6086 279
rect 3744 -217 3753 -146
rect 3824 -217 3833 -146
rect 3744 -226 3833 -217
rect 3556 -306 3646 -295
rect 3556 -374 3567 -306
rect 3635 -374 3646 -306
rect 3556 -385 3646 -374
rect 5287 -893 5571 -879
rect 5287 -1002 5303 -893
rect 5553 -1002 5571 -893
rect 3292 -1058 3576 -1053
rect 3292 -1189 3298 -1058
rect 3565 -1189 3576 -1058
rect -4155 -3444 -3941 -2876
rect -3373 -3444 1204 -2876
rect 3292 -3006 3576 -1189
rect 5287 -2426 5571 -1002
rect 3976 -2482 4399 -2470
rect 3976 -2882 3988 -2482
rect 4388 -2882 4399 -2482
rect 5287 -2716 5571 -2710
rect 5980 -1053 6086 177
rect 6255 162 6261 346
rect 6313 162 6323 346
rect 8668 291 8773 969
rect 12540 831 12928 983
rect 12540 739 12686 831
rect 12778 739 12928 831
rect 12540 586 12928 739
rect 8943 346 9011 353
rect 8668 279 8774 291
rect 6255 -295 6323 162
rect 6432 257 6521 263
rect 6432 179 6438 257
rect 6513 179 6521 257
rect 6432 -146 6521 179
rect 8669 177 8674 279
rect 8768 177 8774 279
rect 6432 -217 6441 -146
rect 6512 -217 6521 -146
rect 6432 -226 6521 -217
rect 6244 -306 6334 -295
rect 6244 -374 6255 -306
rect 6323 -374 6334 -306
rect 6244 -385 6334 -374
rect 7975 -903 8259 -879
rect 7975 -1007 8001 -903
rect 8222 -1007 8259 -903
rect 5980 -1073 6264 -1053
rect 5980 -1189 5986 -1073
rect 6253 -1189 6264 -1073
rect 3976 -2893 4399 -2882
rect 5980 -2725 6264 -1189
rect 7975 -2426 8259 -1007
rect 7975 -2716 8259 -2710
rect 8668 -1053 8774 177
rect 8943 162 8949 346
rect 9001 162 9011 346
rect 11356 279 11462 291
rect 8943 -295 9011 162
rect 9120 257 9209 263
rect 9120 179 9126 257
rect 9201 179 9209 257
rect 9120 -146 9209 179
rect 9120 -217 9129 -146
rect 9200 -217 9209 -146
rect 9120 -226 9209 -217
rect 11356 177 11362 279
rect 11456 177 11462 279
rect 8932 -306 9022 -295
rect 8932 -374 8943 -306
rect 9011 -374 9022 -306
rect 8932 -385 9022 -374
rect 10663 -903 10947 -879
rect 10663 -1006 10686 -903
rect 10902 -1006 10947 -903
rect 8668 -1072 8952 -1053
rect 8668 -1159 8692 -1072
rect 8926 -1159 8952 -1072
rect 3292 -3296 3576 -3290
rect -4155 -3608 -3272 -3444
rect 636 -3523 1204 -3444
rect 636 -3621 3374 -3523
rect 636 -3656 1974 -3621
rect 636 -3729 642 -3656
rect 1967 -3729 1974 -3656
rect 636 -3735 1974 -3729
rect 636 -3875 694 -3735
rect 636 -4862 639 -3875
rect 692 -4862 694 -3875
rect 636 -4868 694 -4862
rect 764 -3875 822 -3868
rect 764 -4862 767 -3875
rect 820 -4862 822 -3875
rect 360 -4903 432 -4898
rect 360 -4909 682 -4903
rect 360 -4912 620 -4909
rect 360 -4968 368 -4912
rect 424 -4965 620 -4912
rect 676 -4965 682 -4909
rect 424 -4968 682 -4965
rect 360 -4971 682 -4968
rect 360 -4974 432 -4971
rect -1245 -5020 -785 -4990
rect 764 -5020 822 -4862
rect 892 -3875 950 -3735
rect 892 -4862 895 -3875
rect 948 -4862 950 -3875
rect 892 -4868 950 -4862
rect 1020 -3875 1078 -3868
rect 1020 -4862 1023 -3875
rect 1076 -4862 1078 -3875
rect 1020 -5020 1078 -4862
rect 1148 -3875 1206 -3735
rect 1148 -4862 1151 -3875
rect 1204 -4862 1206 -3875
rect 1148 -4868 1206 -4862
rect 1276 -3875 1334 -3868
rect 1276 -4862 1279 -3875
rect 1332 -4862 1334 -3875
rect 1276 -5020 1334 -4862
rect 1404 -3875 1462 -3735
rect 1404 -4862 1407 -3875
rect 1460 -4862 1462 -3875
rect 1404 -4868 1462 -4862
rect 1532 -3875 1590 -3868
rect 1532 -4862 1535 -3875
rect 1588 -4862 1590 -3875
rect 1532 -5020 1590 -4862
rect 1660 -3875 1718 -3735
rect 1660 -4862 1663 -3875
rect 1716 -4862 1718 -3875
rect 1660 -4868 1718 -4862
rect 1788 -3875 1846 -3868
rect 1788 -4862 1791 -3875
rect 1844 -4862 1846 -3875
rect 1788 -5020 1846 -4862
rect 1916 -3875 1974 -3735
rect 1916 -4862 1919 -3875
rect 1972 -4862 1974 -3875
rect 1916 -4868 1974 -4862
rect 2348 -4473 2414 -3621
rect 2540 -4473 2606 -3621
rect 2732 -4473 2798 -3621
rect 2924 -4473 2990 -3621
rect 3116 -4473 3182 -3621
rect 3308 -4473 3374 -3621
rect 3541 -3888 3646 -3863
rect 3541 -3944 3563 -3888
rect 3619 -3944 3646 -3888
rect 3541 -3961 3646 -3944
rect 2348 -4867 2354 -4473
rect 2408 -4867 2414 -4473
rect 2348 -4873 2414 -4867
rect 2444 -4867 2450 -4473
rect 2504 -4867 2510 -4473
rect 1904 -4907 2396 -4901
rect 1904 -4909 1911 -4907
rect 1896 -4960 1911 -4909
rect 1983 -4908 2396 -4907
rect 1983 -4960 2338 -4908
rect 1896 -4961 2338 -4960
rect 2390 -4961 2396 -4908
rect 1896 -4965 2396 -4961
rect 2332 -4967 2396 -4965
rect 2444 -5011 2510 -4867
rect 2540 -4867 2546 -4473
rect 2600 -4867 2606 -4473
rect 2540 -4873 2606 -4867
rect 2636 -4867 2642 -4473
rect 2696 -4867 2702 -4473
rect 2636 -5011 2702 -4867
rect 2732 -4867 2738 -4473
rect 2792 -4867 2798 -4473
rect 2732 -4873 2798 -4867
rect 2828 -4867 2834 -4473
rect 2888 -4867 2894 -4473
rect 2828 -5011 2894 -4867
rect 2924 -4867 2930 -4473
rect 2984 -4867 2990 -4473
rect 2924 -4873 2990 -4867
rect 3020 -4867 3026 -4473
rect 3080 -4867 3086 -4473
rect 3020 -5011 3086 -4867
rect 3116 -4867 3122 -4473
rect 3176 -4867 3182 -4473
rect 3116 -4873 3182 -4867
rect 3212 -4867 3218 -4473
rect 3272 -4867 3278 -4473
rect 3212 -5011 3278 -4867
rect 3308 -4867 3314 -4473
rect 3368 -4867 3374 -4473
rect 3308 -4873 3374 -4867
rect 3558 -4901 3628 -3961
rect 3314 -4907 3628 -4901
rect 3314 -4963 3320 -4907
rect 3390 -4963 3628 -4907
rect 3314 -4971 3628 -4963
rect 3988 -5011 4388 -2893
rect 5980 -3015 6264 -3009
rect 8668 -3024 8952 -1159
rect 10663 -2426 10947 -1006
rect 10663 -2716 10947 -2710
rect 11356 -1053 11462 177
rect 16538 -130 17110 1487
rect 19038 720 19500 784
rect 19038 400 19140 720
rect 19460 400 19500 720
rect 19038 337 19500 400
rect 19171 67 19429 337
rect 19160 52 19437 67
rect 19160 -206 19171 52
rect 19429 -206 19437 52
rect 19160 -216 19437 -206
rect 19296 -615 19671 -608
rect 19296 -802 19302 -615
rect 19354 -802 19671 -615
rect 19296 -808 19671 -802
rect 19196 -862 19296 -849
rect 11356 -1078 11640 -1053
rect 11356 -1166 11378 -1078
rect 11608 -1166 11640 -1078
rect 17925 -1110 18390 -929
rect 19196 -933 19206 -862
rect 19286 -933 19296 -862
rect 19196 -943 19296 -933
rect 19208 -1110 19296 -943
rect 8660 -3032 8959 -3024
rect 8660 -3316 8668 -3032
rect 8952 -3316 8959 -3032
rect 8660 -3323 8959 -3316
rect 11356 -3192 11640 -1166
rect 12873 -1149 12943 -1143
rect 12873 -2566 12943 -1219
rect 17925 -1198 18147 -1110
rect 18235 -1198 19296 -1110
rect 17925 -1367 18390 -1198
rect 19208 -1336 19296 -1198
rect 19471 -1065 19671 -808
rect 19471 -1265 41080 -1065
rect 19208 -1347 19308 -1336
rect 19208 -1414 19217 -1347
rect 19298 -1414 19308 -1347
rect 19208 -1425 19308 -1414
rect 19471 -1457 19671 -1265
rect 19308 -1466 19671 -1457
rect 18769 -1483 18951 -1471
rect 18769 -1648 18779 -1483
rect 18944 -1648 18951 -1483
rect 18769 -1654 18951 -1648
rect 19308 -1650 19315 -1466
rect 19367 -1650 19671 -1466
rect 14187 -2043 14277 -1892
rect 14187 -2139 14277 -2133
rect 15150 -2240 15750 -2040
rect 18779 -2240 18944 -1654
rect 19308 -1657 19671 -1650
rect 15150 -2405 18944 -2240
rect 12312 -2572 13512 -2566
rect 12312 -2630 12320 -2572
rect 12736 -2630 13088 -2572
rect 13504 -2630 13512 -2572
rect 12312 -2636 13512 -2630
rect 13842 -2572 14612 -2566
rect 13842 -2630 13850 -2572
rect 14266 -2630 14612 -2572
rect 13842 -2636 14612 -2630
rect 14682 -2636 14691 -2566
rect 11356 -3482 11640 -3476
rect -1245 -5420 -1215 -5020
rect -815 -5420 1846 -5020
rect 2443 -5411 4388 -5011
rect -1245 -5450 -785 -5420
rect 636 -5567 694 -5560
rect 636 -6554 639 -5567
rect 692 -6554 694 -5567
rect 636 -6809 694 -6554
rect 764 -5567 822 -5420
rect 764 -6554 767 -5567
rect 820 -6554 822 -5567
rect 764 -6560 822 -6554
rect 892 -5567 950 -5560
rect 892 -6554 895 -5567
rect 948 -6554 950 -5567
rect 892 -6809 950 -6554
rect 1020 -5567 1078 -5420
rect 1020 -6554 1023 -5567
rect 1076 -6554 1078 -5567
rect 1020 -6560 1078 -6554
rect 1148 -5567 1206 -5560
rect 1148 -6554 1151 -5567
rect 1204 -6554 1206 -5567
rect 1148 -6809 1206 -6554
rect 1276 -5567 1334 -5420
rect 1276 -6554 1279 -5567
rect 1332 -6554 1334 -5567
rect 1276 -6560 1334 -6554
rect 1404 -5567 1462 -5560
rect 1404 -6554 1407 -5567
rect 1460 -6554 1462 -5567
rect 1404 -6809 1462 -6554
rect 1532 -5567 1590 -5420
rect 1532 -6554 1535 -5567
rect 1588 -6554 1590 -5567
rect 1532 -6560 1590 -6554
rect 1660 -5567 1718 -5560
rect 1660 -6554 1663 -5567
rect 1716 -6554 1718 -5567
rect 1660 -6809 1718 -6554
rect 1788 -5567 1846 -5420
rect 2324 -5455 2409 -5454
rect 1902 -5460 2409 -5455
rect 1902 -5461 2331 -5460
rect 1902 -5514 1909 -5461
rect 1981 -5513 2331 -5461
rect 2403 -5513 2409 -5460
rect 1981 -5514 2409 -5513
rect 1902 -5519 2409 -5514
rect 1788 -6554 1791 -5567
rect 1844 -6554 1846 -5567
rect 1788 -6560 1846 -6554
rect 1916 -5567 1974 -5560
rect 1916 -6554 1919 -5567
rect 1972 -6554 1974 -5567
rect 2444 -6351 2508 -5411
rect 2636 -6351 2700 -5411
rect 2828 -6351 2892 -5411
rect 3020 -6351 3084 -5411
rect 3212 -6351 3276 -5411
rect 3312 -5770 3838 -5757
rect 3312 -5776 3683 -5770
rect 3312 -5909 3322 -5776
rect 3374 -5909 3683 -5776
rect 3822 -5909 3838 -5770
rect 3312 -5923 3838 -5909
rect 1916 -6809 1974 -6554
rect -6172 -7150 -5411 -6864
rect -6172 -7536 -6013 -7150
rect -5627 -7536 -5411 -7150
rect -6172 -7739 -5411 -7536
rect 636 -7331 1974 -6809
rect 2348 -6545 2354 -6351
rect 2408 -6545 2414 -6351
rect 2348 -6671 2414 -6545
rect 2444 -6545 2450 -6351
rect 2504 -6545 2510 -6351
rect 2444 -6551 2510 -6545
rect 2540 -6545 2546 -6351
rect 2600 -6545 2606 -6351
rect 2540 -6671 2606 -6545
rect 2636 -6545 2642 -6351
rect 2696 -6545 2702 -6351
rect 2636 -6551 2702 -6545
rect 2732 -6545 2738 -6351
rect 2792 -6545 2798 -6351
rect 2732 -6671 2798 -6545
rect 2828 -6545 2834 -6351
rect 2888 -6545 2894 -6351
rect 2828 -6551 2894 -6545
rect 2924 -6545 2930 -6351
rect 2984 -6545 2990 -6351
rect 2924 -6671 2990 -6545
rect 3020 -6545 3026 -6351
rect 3080 -6545 3086 -6351
rect 3020 -6551 3086 -6545
rect 3116 -6545 3122 -6351
rect 3176 -6545 3182 -6351
rect 3116 -6671 3182 -6545
rect 3212 -6545 3218 -6351
rect 3272 -6545 3278 -6351
rect 3212 -6551 3278 -6545
rect 3308 -6545 3314 -6351
rect 3368 -6398 3374 -6351
rect 15150 -6398 15750 -2405
rect 3368 -6545 15750 -6398
rect 3308 -6671 15750 -6545
rect 2348 -6677 15750 -6671
rect 2348 -6755 2354 -6677
rect 2792 -6755 2930 -6677
rect 3368 -6755 15750 -6677
rect 2348 -6988 15750 -6755
rect 2348 -7150 2391 -6988
rect 3339 -6998 15750 -6988
rect 3339 -7150 3374 -6998
rect 2348 -7176 3374 -7150
rect 636 -7931 40578 -7331
rect 39978 -11865 40578 -7931
rect 40880 -11340 41080 -1265
rect 40880 -11540 42133 -11340
rect 42032 -11849 42133 -11540
rect 41191 -11865 41991 -11859
rect 39978 -11867 41991 -11865
rect 39978 -11921 41203 -11867
rect 41979 -11921 41991 -11867
rect 39978 -11923 41991 -11921
rect 39978 -12181 40578 -11923
rect 41191 -11929 41991 -11923
rect 42032 -11916 42050 -11849
rect 42114 -11916 42133 -11849
rect 42032 -11934 42133 -11916
rect 41191 -12023 41991 -12017
rect 42425 -12023 42537 -12016
rect 41191 -12025 42538 -12023
rect 41191 -12079 41203 -12025
rect 41979 -12036 42538 -12025
rect 41979 -12079 42450 -12036
rect 41191 -12081 42450 -12079
rect 41191 -12087 41991 -12081
rect 42425 -12096 42450 -12081
rect 42510 -12096 42538 -12036
rect 42425 -12114 42538 -12096
rect 41191 -12181 41991 -12175
rect 39978 -12183 41991 -12181
rect 39978 -12237 41203 -12183
rect 41979 -12237 41991 -12183
rect 39978 -12239 41991 -12237
rect 39978 -12497 40578 -12239
rect 41191 -12245 41991 -12239
rect 41191 -12339 41991 -12333
rect 42480 -12339 42538 -12114
rect 41191 -12341 42538 -12339
rect 41191 -12395 41203 -12341
rect 41979 -12395 42538 -12341
rect 41191 -12397 42538 -12395
rect 41191 -12403 41991 -12397
rect 41191 -12497 41991 -12491
rect 39978 -12499 41991 -12497
rect 39978 -12553 41203 -12499
rect 41979 -12553 41991 -12499
rect 39978 -12555 41991 -12553
rect 39978 -12813 40578 -12555
rect 41191 -12561 41991 -12555
rect 41191 -12655 41991 -12649
rect 42480 -12655 42538 -12397
rect 41191 -12657 42538 -12655
rect 41191 -12711 41203 -12657
rect 41979 -12711 42538 -12657
rect 41191 -12713 42538 -12711
rect 41191 -12719 41991 -12713
rect 41191 -12813 41991 -12807
rect 39978 -12815 41991 -12813
rect 39978 -12869 41203 -12815
rect 41979 -12869 41991 -12815
rect 39978 -12871 41991 -12869
rect 39978 -13129 40578 -12871
rect 41191 -12877 41991 -12871
rect 41191 -12971 41991 -12965
rect 42480 -12971 42538 -12713
rect 41191 -12973 42538 -12971
rect 41191 -13027 41203 -12973
rect 41979 -13027 42538 -12973
rect 41191 -13029 42538 -13027
rect 41191 -13035 41991 -13029
rect 41191 -13129 41991 -13123
rect 39978 -13131 41991 -13129
rect 39978 -13185 41203 -13131
rect 41979 -13185 41991 -13131
rect 39978 -13187 41991 -13185
rect 39978 -13445 40578 -13187
rect 41191 -13193 41991 -13187
rect 41191 -13287 41991 -13281
rect 42480 -13287 42538 -13029
rect 41191 -13289 42538 -13287
rect 41191 -13343 41203 -13289
rect 41979 -13343 42538 -13289
rect 41191 -13345 42538 -13343
rect 41191 -13351 41991 -13345
rect 41191 -13445 41991 -13439
rect 39978 -13447 41991 -13445
rect 39978 -13501 41203 -13447
rect 41979 -13501 41991 -13447
rect 39978 -13503 41991 -13501
rect 39978 -13761 40578 -13503
rect 41191 -13509 41991 -13503
rect 41191 -13603 41991 -13597
rect 42480 -13603 42538 -13345
rect 41191 -13605 42538 -13603
rect 41191 -13659 41203 -13605
rect 41979 -13659 42538 -13605
rect 41191 -13661 42538 -13659
rect 41191 -13667 41991 -13661
rect 41191 -13761 41991 -13755
rect 39978 -13763 41991 -13761
rect 39978 -13817 41203 -13763
rect 41979 -13817 41991 -13763
rect 39978 -13819 41991 -13817
rect 39978 -14077 40578 -13819
rect 41191 -13825 41991 -13819
rect 41191 -13919 41991 -13913
rect 42480 -13919 42538 -13661
rect 41191 -13921 42538 -13919
rect 41191 -13975 41203 -13921
rect 41979 -13975 42538 -13921
rect 41191 -13977 42538 -13975
rect 41191 -13983 41991 -13977
rect 41191 -14077 41991 -14071
rect 39978 -14079 41991 -14077
rect 39978 -14133 41203 -14079
rect 41979 -14133 41991 -14079
rect 39978 -14135 41991 -14133
rect 39978 -14393 40578 -14135
rect 41191 -14141 41991 -14135
rect 41191 -14235 41991 -14229
rect 42480 -14235 42538 -13977
rect 41191 -14237 42538 -14235
rect 41191 -14291 41203 -14237
rect 41979 -14291 42538 -14237
rect 41191 -14293 42538 -14291
rect 41191 -14299 41991 -14293
rect 41191 -14393 41991 -14387
rect 39978 -14395 41991 -14393
rect 39978 -14449 41203 -14395
rect 41979 -14449 41991 -14395
rect 39978 -14451 41991 -14449
rect 39978 -14709 40578 -14451
rect 41191 -14457 41991 -14451
rect 41191 -14551 41991 -14545
rect 42480 -14551 42538 -14293
rect 41191 -14553 42538 -14551
rect 41191 -14607 41203 -14553
rect 41979 -14607 42538 -14553
rect 41191 -14609 42538 -14607
rect 41191 -14615 41991 -14609
rect 41191 -14709 41991 -14703
rect 39978 -14711 41991 -14709
rect 39978 -14765 41203 -14711
rect 41979 -14765 41991 -14711
rect 39978 -14767 41991 -14765
rect 39978 -15025 40578 -14767
rect 41191 -14773 41991 -14767
rect 41191 -14867 41991 -14861
rect 42480 -14867 42538 -14609
rect 41191 -14869 42538 -14867
rect 41191 -14923 41203 -14869
rect 41979 -14923 42538 -14869
rect 41191 -14925 42538 -14923
rect 41191 -14931 41991 -14925
rect 41191 -15025 41991 -15019
rect 39978 -15027 41991 -15025
rect 39978 -15081 41203 -15027
rect 41979 -15081 41991 -15027
rect 39978 -15083 41991 -15081
rect 39978 -15341 40578 -15083
rect 41191 -15089 41991 -15083
rect 41191 -15183 41991 -15177
rect 42480 -15183 42538 -14925
rect 41191 -15185 42538 -15183
rect 41191 -15239 41203 -15185
rect 41979 -15239 42538 -15185
rect 41191 -15241 42538 -15239
rect 41191 -15247 41991 -15241
rect 41191 -15341 41991 -15335
rect 39978 -15343 41991 -15341
rect 39978 -15397 41203 -15343
rect 41979 -15397 41991 -15343
rect 39978 -15399 41991 -15397
rect 39978 -15657 40578 -15399
rect 41191 -15405 41991 -15399
rect 41191 -15499 41991 -15493
rect 42480 -15499 42538 -15241
rect 41191 -15501 42538 -15499
rect 41191 -15555 41203 -15501
rect 41979 -15555 42538 -15501
rect 41191 -15557 42538 -15555
rect 41191 -15563 41991 -15557
rect 41191 -15657 41991 -15651
rect 39978 -15659 41991 -15657
rect 39978 -15713 41203 -15659
rect 41979 -15713 41991 -15659
rect 39978 -15715 41991 -15713
rect 39978 -15973 40578 -15715
rect 41191 -15721 41991 -15715
rect 41191 -15815 41991 -15809
rect 42480 -15815 42538 -15557
rect 41191 -15817 42538 -15815
rect 41191 -15871 41203 -15817
rect 41979 -15871 42538 -15817
rect 41191 -15873 42538 -15871
rect 41191 -15879 41991 -15873
rect 41191 -15973 41991 -15967
rect 39978 -15975 41991 -15973
rect 39978 -16029 41203 -15975
rect 41979 -16029 41991 -15975
rect 39978 -16031 41991 -16029
rect 39978 -16289 40578 -16031
rect 41191 -16037 41991 -16031
rect 41191 -16131 41991 -16125
rect 42480 -16131 42538 -15873
rect 41191 -16133 42538 -16131
rect 41191 -16187 41203 -16133
rect 41979 -16187 42538 -16133
rect 41191 -16189 42538 -16187
rect 41191 -16195 41991 -16189
rect 41191 -16289 41991 -16283
rect 39978 -16291 41991 -16289
rect 39978 -16345 41203 -16291
rect 41979 -16345 41991 -16291
rect 39978 -16347 41991 -16345
rect 4080 -16482 4399 -16470
rect -4155 -16876 -3272 -16759
rect -4155 -17444 -3941 -16876
rect -3373 -16878 -1892 -16876
rect -3373 -17444 1204 -16878
rect -4155 -17608 -3272 -17444
rect 636 -17523 1204 -17444
rect 3988 -16882 4080 -16698
rect 4388 -16882 4399 -16482
rect 3988 -16893 4399 -16882
rect 39978 -16605 40578 -16347
rect 41191 -16353 41991 -16347
rect 41191 -16447 41991 -16441
rect 42480 -16447 42538 -16189
rect 41191 -16449 42538 -16447
rect 41191 -16503 41203 -16449
rect 41979 -16503 42538 -16449
rect 41191 -16505 42538 -16503
rect 41191 -16511 41991 -16505
rect 41191 -16605 41991 -16599
rect 39978 -16607 41991 -16605
rect 39978 -16661 41203 -16607
rect 41979 -16661 41991 -16607
rect 39978 -16663 41991 -16661
rect 636 -17621 3374 -17523
rect 636 -17656 1974 -17621
rect 636 -17729 642 -17656
rect 1967 -17729 1974 -17656
rect 636 -17735 1974 -17729
rect 636 -17875 694 -17735
rect 636 -18862 639 -17875
rect 692 -18862 694 -17875
rect 636 -18868 694 -18862
rect 764 -17875 822 -17868
rect 764 -18862 767 -17875
rect 820 -18862 822 -17875
rect 360 -18903 432 -18898
rect 360 -18909 682 -18903
rect 360 -18912 620 -18909
rect 360 -18968 368 -18912
rect 424 -18965 620 -18912
rect 676 -18965 682 -18909
rect 424 -18968 682 -18965
rect 360 -18971 682 -18968
rect 360 -18974 432 -18971
rect -1245 -19020 -785 -18990
rect 764 -19020 822 -18862
rect 892 -17875 950 -17735
rect 892 -18862 895 -17875
rect 948 -18862 950 -17875
rect 892 -18868 950 -18862
rect 1020 -17875 1078 -17868
rect 1020 -18862 1023 -17875
rect 1076 -18862 1078 -17875
rect 1020 -19020 1078 -18862
rect 1148 -17875 1206 -17735
rect 1148 -18862 1151 -17875
rect 1204 -18862 1206 -17875
rect 1148 -18868 1206 -18862
rect 1276 -17875 1334 -17868
rect 1276 -18862 1279 -17875
rect 1332 -18862 1334 -17875
rect 1276 -19020 1334 -18862
rect 1404 -17875 1462 -17735
rect 1404 -18862 1407 -17875
rect 1460 -18862 1462 -17875
rect 1404 -18868 1462 -18862
rect 1532 -17875 1590 -17868
rect 1532 -18862 1535 -17875
rect 1588 -18862 1590 -17875
rect 1532 -19020 1590 -18862
rect 1660 -17875 1718 -17735
rect 1660 -18862 1663 -17875
rect 1716 -18862 1718 -17875
rect 1660 -18868 1718 -18862
rect 1788 -17875 1846 -17868
rect 1788 -18862 1791 -17875
rect 1844 -18862 1846 -17875
rect 1788 -19020 1846 -18862
rect 1916 -17875 1974 -17735
rect 1916 -18862 1919 -17875
rect 1972 -18862 1974 -17875
rect 1916 -18868 1974 -18862
rect 2348 -18473 2414 -17621
rect 2540 -18473 2606 -17621
rect 2732 -18473 2798 -17621
rect 2924 -18473 2990 -17621
rect 3116 -18473 3182 -17621
rect 3308 -18473 3374 -17621
rect 3541 -17888 3646 -17863
rect 3541 -17944 3563 -17888
rect 3619 -17944 3646 -17888
rect 3541 -17961 3646 -17944
rect 2348 -18867 2354 -18473
rect 2408 -18867 2414 -18473
rect 2348 -18873 2414 -18867
rect 2444 -18867 2450 -18473
rect 2504 -18867 2510 -18473
rect 1904 -18907 2396 -18901
rect 1904 -18909 1911 -18907
rect 1896 -18960 1911 -18909
rect 1983 -18908 2396 -18907
rect 1983 -18960 2338 -18908
rect 1896 -18961 2338 -18960
rect 2390 -18961 2396 -18908
rect 1896 -18965 2396 -18961
rect 2332 -18967 2396 -18965
rect 2444 -19011 2510 -18867
rect 2540 -18867 2546 -18473
rect 2600 -18867 2606 -18473
rect 2540 -18873 2606 -18867
rect 2636 -18867 2642 -18473
rect 2696 -18867 2702 -18473
rect 2636 -19011 2702 -18867
rect 2732 -18867 2738 -18473
rect 2792 -18867 2798 -18473
rect 2732 -18873 2798 -18867
rect 2828 -18867 2834 -18473
rect 2888 -18867 2894 -18473
rect 2828 -19011 2894 -18867
rect 2924 -18867 2930 -18473
rect 2984 -18867 2990 -18473
rect 2924 -18873 2990 -18867
rect 3020 -18867 3026 -18473
rect 3080 -18867 3086 -18473
rect 3020 -19011 3086 -18867
rect 3116 -18867 3122 -18473
rect 3176 -18867 3182 -18473
rect 3116 -18873 3182 -18867
rect 3212 -18867 3218 -18473
rect 3272 -18867 3278 -18473
rect 3212 -19011 3278 -18867
rect 3308 -18867 3314 -18473
rect 3368 -18867 3374 -18473
rect 3308 -18873 3374 -18867
rect 3558 -18901 3628 -17961
rect 3314 -18907 3628 -18901
rect 3314 -18963 3320 -18907
rect 3390 -18963 3628 -18907
rect 3314 -18971 3628 -18963
rect 3988 -19011 4388 -16893
rect -1245 -19420 -1215 -19020
rect -815 -19420 1846 -19020
rect 2443 -19411 4388 -19011
rect 39978 -16921 40578 -16663
rect 41191 -16669 41991 -16663
rect 41191 -16763 41991 -16757
rect 42480 -16763 42538 -16505
rect 41191 -16765 42538 -16763
rect 41191 -16819 41203 -16765
rect 41979 -16819 42538 -16765
rect 41191 -16821 42538 -16819
rect 41191 -16827 41991 -16821
rect 41191 -16921 41991 -16915
rect 39978 -16923 41991 -16921
rect 39978 -16977 41203 -16923
rect 41979 -16977 41991 -16923
rect 39978 -16979 41991 -16977
rect 39978 -17237 40578 -16979
rect 41191 -16985 41991 -16979
rect 41191 -17079 41991 -17073
rect 42480 -17079 42538 -16821
rect 41191 -17081 42538 -17079
rect 41191 -17135 41203 -17081
rect 41979 -17135 42538 -17081
rect 41191 -17137 42538 -17135
rect 41191 -17143 41991 -17137
rect 41191 -17237 41991 -17231
rect 39978 -17239 41991 -17237
rect 39978 -17293 41203 -17239
rect 41979 -17293 41991 -17239
rect 39978 -17295 41991 -17293
rect 39978 -17553 40578 -17295
rect 41191 -17301 41991 -17295
rect 41191 -17395 41991 -17389
rect 42480 -17395 42538 -17137
rect 41191 -17397 42538 -17395
rect 41191 -17451 41203 -17397
rect 41979 -17451 42538 -17397
rect 41191 -17453 42538 -17451
rect 41191 -17459 41991 -17453
rect 41191 -17553 41991 -17547
rect 39978 -17555 41991 -17553
rect 39978 -17609 41203 -17555
rect 41979 -17609 41991 -17555
rect 39978 -17611 41991 -17609
rect 39978 -17869 40578 -17611
rect 41191 -17617 41991 -17611
rect 41191 -17711 41991 -17705
rect 42480 -17711 42538 -17453
rect 41191 -17713 42538 -17711
rect 41191 -17767 41203 -17713
rect 41979 -17767 42538 -17713
rect 41191 -17769 42538 -17767
rect 41191 -17775 41991 -17769
rect 41191 -17869 41991 -17863
rect 39978 -17871 41991 -17869
rect 39978 -17925 41203 -17871
rect 41979 -17925 41991 -17871
rect 39978 -17927 41991 -17925
rect 39978 -18185 40578 -17927
rect 41191 -17933 41991 -17927
rect 41191 -18027 41991 -18021
rect 42480 -18027 42538 -17769
rect 41191 -18029 42538 -18027
rect 41191 -18083 41203 -18029
rect 41979 -18083 42538 -18029
rect 41191 -18085 42538 -18083
rect 41191 -18091 41991 -18085
rect 41191 -18185 41991 -18179
rect 39978 -18187 41991 -18185
rect 39978 -18241 41203 -18187
rect 41979 -18241 41991 -18187
rect 39978 -18243 41991 -18241
rect 39978 -18501 40578 -18243
rect 41191 -18249 41991 -18243
rect 41191 -18343 41991 -18337
rect 42480 -18343 42538 -18085
rect 41191 -18345 42538 -18343
rect 41191 -18399 41203 -18345
rect 41979 -18399 42538 -18345
rect 41191 -18401 42538 -18399
rect 41191 -18407 41991 -18401
rect 41191 -18501 41991 -18495
rect 39978 -18503 41991 -18501
rect 39978 -18557 41203 -18503
rect 41979 -18557 41991 -18503
rect 39978 -18559 41991 -18557
rect 39978 -18817 40578 -18559
rect 41191 -18565 41991 -18559
rect 41191 -18659 41991 -18653
rect 42480 -18659 42538 -18401
rect 41191 -18661 42538 -18659
rect 41191 -18715 41203 -18661
rect 41979 -18715 42538 -18661
rect 41191 -18717 42538 -18715
rect 41191 -18723 41991 -18717
rect 41191 -18817 41991 -18811
rect 39978 -18819 41991 -18817
rect 39978 -18873 41203 -18819
rect 41979 -18873 41991 -18819
rect 39978 -18875 41991 -18873
rect 39978 -19133 40578 -18875
rect 41191 -18881 41991 -18875
rect 41191 -18975 41991 -18969
rect 42480 -18975 42538 -18717
rect 41191 -18977 42538 -18975
rect 41191 -19031 41203 -18977
rect 41979 -19031 42538 -18977
rect 41191 -19033 42538 -19031
rect 41191 -19039 41991 -19033
rect 41191 -19133 41991 -19127
rect 39978 -19135 41991 -19133
rect 39978 -19189 41203 -19135
rect 41979 -19189 41991 -19135
rect 39978 -19191 41991 -19189
rect -1245 -19450 -785 -19420
rect 636 -19567 694 -19560
rect 636 -20554 639 -19567
rect 692 -20554 694 -19567
rect 636 -20809 694 -20554
rect 764 -19567 822 -19420
rect 764 -20554 767 -19567
rect 820 -20554 822 -19567
rect 764 -20560 822 -20554
rect 892 -19567 950 -19560
rect 892 -20554 895 -19567
rect 948 -20554 950 -19567
rect 892 -20809 950 -20554
rect 1020 -19567 1078 -19420
rect 1020 -20554 1023 -19567
rect 1076 -20554 1078 -19567
rect 1020 -20560 1078 -20554
rect 1148 -19567 1206 -19560
rect 1148 -20554 1151 -19567
rect 1204 -20554 1206 -19567
rect 1148 -20809 1206 -20554
rect 1276 -19567 1334 -19420
rect 1276 -20554 1279 -19567
rect 1332 -20554 1334 -19567
rect 1276 -20560 1334 -20554
rect 1404 -19567 1462 -19560
rect 1404 -20554 1407 -19567
rect 1460 -20554 1462 -19567
rect 1404 -20809 1462 -20554
rect 1532 -19567 1590 -19420
rect 1532 -20554 1535 -19567
rect 1588 -20554 1590 -19567
rect 1532 -20560 1590 -20554
rect 1660 -19567 1718 -19560
rect 1660 -20554 1663 -19567
rect 1716 -20554 1718 -19567
rect 1660 -20809 1718 -20554
rect 1788 -19567 1846 -19420
rect 2324 -19455 2409 -19454
rect 1902 -19460 2409 -19455
rect 1902 -19461 2331 -19460
rect 1902 -19514 1909 -19461
rect 1981 -19513 2331 -19461
rect 2403 -19513 2409 -19460
rect 1981 -19514 2409 -19513
rect 1902 -19519 2409 -19514
rect 1788 -20554 1791 -19567
rect 1844 -20554 1846 -19567
rect 1788 -20560 1846 -20554
rect 1916 -19567 1974 -19560
rect 1916 -20554 1919 -19567
rect 1972 -20554 1974 -19567
rect 2444 -20351 2508 -19411
rect 2636 -20351 2700 -19411
rect 2828 -20351 2892 -19411
rect 3020 -20351 3084 -19411
rect 3212 -20351 3276 -19411
rect 39978 -19449 40578 -19191
rect 41191 -19197 41991 -19191
rect 41191 -19291 41991 -19285
rect 42480 -19291 42538 -19033
rect 41191 -19293 42538 -19291
rect 41191 -19347 41203 -19293
rect 41979 -19347 42538 -19293
rect 41191 -19349 42538 -19347
rect 41191 -19355 41991 -19349
rect 41191 -19449 41991 -19443
rect 39978 -19451 41991 -19449
rect 39978 -19505 41203 -19451
rect 41979 -19505 41991 -19451
rect 39978 -19507 41991 -19505
rect 3312 -19770 3838 -19757
rect 3312 -19776 3683 -19770
rect 3312 -19909 3322 -19776
rect 3374 -19909 3683 -19776
rect 3822 -19909 3838 -19770
rect 3312 -19923 3838 -19909
rect 39978 -19765 40578 -19507
rect 41191 -19513 41991 -19507
rect 41191 -19607 41991 -19601
rect 42480 -19607 42538 -19349
rect 41191 -19609 42538 -19607
rect 41191 -19663 41203 -19609
rect 41979 -19663 42538 -19609
rect 41191 -19665 42538 -19663
rect 41191 -19671 41991 -19665
rect 41191 -19765 41991 -19759
rect 39978 -19767 41991 -19765
rect 39978 -19821 41203 -19767
rect 41979 -19821 41991 -19767
rect 39978 -19823 41991 -19821
rect 39978 -20081 40578 -19823
rect 41191 -19829 41991 -19823
rect 41191 -19923 41991 -19917
rect 42480 -19923 42538 -19665
rect 41191 -19925 42538 -19923
rect 41191 -19979 41203 -19925
rect 41979 -19979 42538 -19925
rect 41191 -19981 42538 -19979
rect 41191 -19987 41991 -19981
rect 41191 -20081 41991 -20075
rect 39978 -20083 41991 -20081
rect 39978 -20137 41203 -20083
rect 41979 -20137 41991 -20083
rect 39978 -20139 41991 -20137
rect 1916 -20809 1974 -20554
rect -6172 -21150 -5411 -20864
rect -6172 -21536 -6013 -21150
rect -5627 -21536 -5411 -21150
rect -6172 -21739 -5411 -21536
rect 636 -21331 1974 -20809
rect 2348 -20545 2354 -20351
rect 2408 -20545 2414 -20351
rect 2348 -20671 2414 -20545
rect 2444 -20545 2450 -20351
rect 2504 -20545 2510 -20351
rect 2444 -20551 2510 -20545
rect 2540 -20545 2546 -20351
rect 2600 -20545 2606 -20351
rect 2540 -20671 2606 -20545
rect 2636 -20545 2642 -20351
rect 2696 -20545 2702 -20351
rect 2636 -20551 2702 -20545
rect 2732 -20545 2738 -20351
rect 2792 -20545 2798 -20351
rect 2732 -20671 2798 -20545
rect 2828 -20545 2834 -20351
rect 2888 -20545 2894 -20351
rect 2828 -20551 2894 -20545
rect 2924 -20545 2930 -20351
rect 2984 -20545 2990 -20351
rect 2924 -20671 2990 -20545
rect 3020 -20545 3026 -20351
rect 3080 -20545 3086 -20351
rect 3020 -20551 3086 -20545
rect 3116 -20545 3122 -20351
rect 3176 -20545 3182 -20351
rect 3116 -20671 3182 -20545
rect 3212 -20545 3218 -20351
rect 3272 -20545 3278 -20351
rect 3212 -20551 3278 -20545
rect 3308 -20545 3314 -20351
rect 3368 -20545 3374 -20351
rect 3308 -20671 3374 -20545
rect 2348 -20677 3374 -20671
rect 2348 -20755 2354 -20677
rect 2792 -20755 2930 -20677
rect 3368 -20755 3374 -20677
rect 2348 -20988 3374 -20755
rect 2348 -21150 2391 -20988
rect 3339 -21150 3374 -20988
rect 2348 -21176 3374 -21150
rect 39978 -20397 40578 -20139
rect 41191 -20145 41991 -20139
rect 41191 -20239 41991 -20233
rect 42480 -20239 42538 -19981
rect 41191 -20241 42538 -20239
rect 41191 -20295 41203 -20241
rect 41979 -20295 42538 -20241
rect 41191 -20297 42538 -20295
rect 41191 -20303 41991 -20297
rect 41191 -20397 41991 -20391
rect 39978 -20399 41991 -20397
rect 39978 -20453 41203 -20399
rect 41979 -20453 41991 -20399
rect 39978 -20455 41991 -20453
rect 39978 -20713 40578 -20455
rect 41191 -20461 41991 -20455
rect 41191 -20555 41991 -20549
rect 42480 -20555 42538 -20297
rect 41191 -20557 42538 -20555
rect 41191 -20611 41203 -20557
rect 41979 -20611 42538 -20557
rect 41191 -20613 42538 -20611
rect 41191 -20619 41991 -20613
rect 41191 -20713 41991 -20707
rect 39978 -20715 41991 -20713
rect 39978 -20769 41203 -20715
rect 41979 -20769 41991 -20715
rect 39978 -20771 41991 -20769
rect 39978 -21029 40578 -20771
rect 41191 -20777 41991 -20771
rect 41191 -20871 41991 -20865
rect 42480 -20871 42538 -20613
rect 41191 -20873 42538 -20871
rect 41191 -20927 41203 -20873
rect 41979 -20927 42538 -20873
rect 41191 -20929 42538 -20927
rect 41191 -20935 41991 -20929
rect 41191 -21029 41991 -21023
rect 39978 -21031 41991 -21029
rect 39978 -21085 41203 -21031
rect 41979 -21085 41991 -21031
rect 39978 -21087 41991 -21085
rect 39978 -21331 40578 -21087
rect 41191 -21093 41991 -21087
rect 41191 -21187 41991 -21181
rect 42480 -21187 42538 -20929
rect 41191 -21189 42538 -21187
rect 41191 -21243 41203 -21189
rect 41979 -21243 42538 -21189
rect 41191 -21245 42538 -21243
rect 41191 -21251 41991 -21245
rect 636 -21345 40578 -21331
rect 41191 -21345 41991 -21339
rect 636 -21347 41991 -21345
rect 636 -21401 41203 -21347
rect 41979 -21401 41991 -21347
rect 636 -21403 41991 -21401
rect 636 -21661 40578 -21403
rect 41191 -21409 41991 -21403
rect 41191 -21503 41991 -21497
rect 42480 -21503 42538 -21245
rect 41191 -21505 42538 -21503
rect 41191 -21559 41203 -21505
rect 41979 -21559 42538 -21505
rect 41191 -21561 42538 -21559
rect 41191 -21567 41991 -21561
rect 41191 -21661 41991 -21655
rect 636 -21663 41991 -21661
rect 636 -21717 41203 -21663
rect 41979 -21717 41991 -21663
rect 636 -21719 41991 -21717
rect 636 -21931 40578 -21719
rect 41191 -21725 41991 -21719
rect 41191 -21819 41991 -21813
rect 42480 -21819 42538 -21561
rect 41191 -21821 42538 -21819
rect 41191 -21875 41203 -21821
rect 41979 -21875 42538 -21821
rect 41191 -21877 42538 -21875
rect 41191 -21883 41991 -21877
rect 39978 -21977 40578 -21931
rect 41191 -21977 41991 -21971
rect 39978 -21979 41991 -21977
rect 39978 -22033 41203 -21979
rect 41979 -22033 41991 -21979
rect 39978 -22035 41991 -22033
rect 39978 -22293 40578 -22035
rect 41191 -22041 41991 -22035
rect 41191 -22135 41991 -22129
rect 42480 -22135 42538 -21877
rect 41191 -22137 42538 -22135
rect 41191 -22191 41203 -22137
rect 41979 -22191 42538 -22137
rect 41191 -22193 42538 -22191
rect 41191 -22199 41991 -22193
rect 41191 -22293 41991 -22287
rect 39978 -22295 41991 -22293
rect 39978 -22349 41203 -22295
rect 41979 -22349 41991 -22295
rect 39978 -22351 41991 -22349
rect 39978 -22609 40578 -22351
rect 41191 -22357 41991 -22351
rect 41191 -22451 41991 -22445
rect 42480 -22451 42538 -22193
rect 41191 -22453 42538 -22451
rect 41191 -22507 41203 -22453
rect 41979 -22507 42538 -22453
rect 41191 -22509 42538 -22507
rect 41191 -22515 41991 -22509
rect 41191 -22609 41991 -22603
rect 39978 -22611 41991 -22609
rect 39978 -22665 41203 -22611
rect 41979 -22665 41991 -22611
rect 39978 -22667 41991 -22665
rect 39978 -22925 40578 -22667
rect 41191 -22673 41991 -22667
rect 41191 -22767 41991 -22761
rect 42480 -22767 42538 -22509
rect 41191 -22769 42538 -22767
rect 41191 -22823 41203 -22769
rect 41979 -22823 42538 -22769
rect 41191 -22825 42538 -22823
rect 41191 -22831 41991 -22825
rect 41191 -22925 41991 -22919
rect 39978 -22927 41991 -22925
rect 39978 -22981 41203 -22927
rect 41979 -22981 41991 -22927
rect 39978 -22983 41991 -22981
rect 39978 -23241 40578 -22983
rect 41191 -22989 41991 -22983
rect 41191 -23083 41991 -23077
rect 42480 -23083 42538 -22825
rect 41191 -23085 42538 -23083
rect 41191 -23139 41203 -23085
rect 41979 -23139 42538 -23085
rect 41191 -23141 42538 -23139
rect 41191 -23147 41991 -23141
rect 41191 -23241 41991 -23235
rect 39978 -23243 41991 -23241
rect 39978 -23297 41203 -23243
rect 41979 -23297 41991 -23243
rect 39978 -23299 41991 -23297
rect 39978 -23557 40578 -23299
rect 41191 -23305 41991 -23299
rect 41191 -23399 41991 -23393
rect 42480 -23399 42538 -23141
rect 41191 -23401 42538 -23399
rect 41191 -23455 41203 -23401
rect 41979 -23455 42538 -23401
rect 41191 -23457 42538 -23455
rect 41191 -23463 41991 -23457
rect 41191 -23557 41991 -23551
rect 39978 -23559 41991 -23557
rect 39978 -23613 41203 -23559
rect 41979 -23613 41991 -23559
rect 39978 -23615 41991 -23613
rect 39978 -23873 40578 -23615
rect 41191 -23621 41991 -23615
rect 41191 -23715 41991 -23709
rect 42480 -23715 42538 -23457
rect 41191 -23717 42538 -23715
rect 41191 -23771 41203 -23717
rect 41979 -23771 42538 -23717
rect 41191 -23773 42538 -23771
rect 41191 -23779 41991 -23773
rect 41191 -23873 41991 -23867
rect 39978 -23875 41991 -23873
rect 39978 -23929 41203 -23875
rect 41979 -23929 41991 -23875
rect 39978 -23931 41991 -23929
rect 39978 -24189 40578 -23931
rect 41191 -23937 41991 -23931
rect 41191 -24031 41991 -24025
rect 42480 -24031 42538 -23773
rect 41191 -24033 42538 -24031
rect 41191 -24087 41203 -24033
rect 41979 -24087 42538 -24033
rect 41191 -24089 42538 -24087
rect 41191 -24095 41991 -24089
rect 41191 -24189 41991 -24183
rect 39978 -24191 41991 -24189
rect 39978 -24245 41203 -24191
rect 41979 -24245 41991 -24191
rect 39978 -24247 41991 -24245
rect 39978 -24505 40578 -24247
rect 41191 -24253 41991 -24247
rect 41191 -24347 41991 -24341
rect 42480 -24347 42538 -24089
rect 41191 -24349 42538 -24347
rect 41191 -24403 41203 -24349
rect 41979 -24403 42538 -24349
rect 41191 -24405 42538 -24403
rect 41191 -24411 41991 -24405
rect 41191 -24505 41991 -24499
rect 39978 -24507 41991 -24505
rect 39978 -24561 41203 -24507
rect 41979 -24561 41991 -24507
rect 39978 -24563 41991 -24561
rect 39978 -25910 40578 -24563
rect 41191 -24569 41991 -24563
rect 41107 -25440 41349 -25417
rect 41107 -25445 42217 -25440
rect 41107 -25633 41132 -25445
rect 41320 -25633 42217 -25445
rect 41107 -25638 42217 -25633
rect 41107 -25654 41349 -25638
rect 41174 -25910 41974 -25905
rect 39978 -25912 41974 -25910
rect 39978 -25966 41186 -25912
rect 41962 -25966 41974 -25912
rect 42019 -25938 42217 -25638
rect 39978 -25968 41974 -25966
rect 39978 -26226 40578 -25968
rect 41174 -25973 41974 -25968
rect 42006 -25946 42217 -25938
rect 42006 -26014 42014 -25946
rect 42098 -25995 42217 -25946
rect 42098 -26014 42105 -25995
rect 42006 -26023 42105 -26014
rect 41042 -26056 41139 -26047
rect 41042 -26151 41053 -26056
rect 41128 -26151 41139 -26056
rect 41174 -26068 41974 -26063
rect 42480 -26068 42538 -24405
rect 41174 -26070 42538 -26068
rect 41174 -26124 41186 -26070
rect 41962 -26124 42538 -26070
rect 41174 -26126 42538 -26124
rect 41174 -26131 41974 -26126
rect 41042 -26159 41139 -26151
rect 41174 -26226 41974 -26221
rect 39978 -26228 41974 -26226
rect 39978 -26282 41186 -26228
rect 41962 -26282 41974 -26228
rect 39978 -26284 41974 -26282
rect 39978 -26542 40578 -26284
rect 41174 -26289 41974 -26284
rect 41174 -26384 41974 -26379
rect 42480 -26384 42538 -26126
rect 41174 -26386 42538 -26384
rect 41174 -26440 41186 -26386
rect 41962 -26440 42538 -26386
rect 41174 -26442 42538 -26440
rect 41174 -26447 41974 -26442
rect 41174 -26542 41974 -26537
rect 39978 -26544 41974 -26542
rect 39978 -26598 41186 -26544
rect 41962 -26598 41974 -26544
rect 39978 -26600 41974 -26598
rect 39978 -26858 40578 -26600
rect 41174 -26605 41974 -26600
rect 41174 -26700 41974 -26695
rect 42480 -26700 42538 -26442
rect 41174 -26702 42538 -26700
rect 41174 -26756 41186 -26702
rect 41962 -26756 42538 -26702
rect 41174 -26758 42538 -26756
rect 41174 -26763 41974 -26758
rect 41174 -26858 41974 -26853
rect 39978 -26860 41974 -26858
rect 39978 -26914 41186 -26860
rect 41962 -26914 41974 -26860
rect 39978 -26916 41974 -26914
rect 39978 -27174 40578 -26916
rect 41174 -26921 41974 -26916
rect 41174 -27016 41974 -27011
rect 42480 -27016 42538 -26758
rect 41174 -27018 42538 -27016
rect 41174 -27072 41186 -27018
rect 41962 -27072 42538 -27018
rect 41174 -27074 42538 -27072
rect 41174 -27079 41974 -27074
rect 41174 -27174 41974 -27169
rect 39978 -27176 41974 -27174
rect 39978 -27230 41186 -27176
rect 41962 -27230 41974 -27176
rect 39978 -27232 41974 -27230
rect 39978 -27490 40578 -27232
rect 41174 -27237 41974 -27232
rect 41174 -27332 41974 -27327
rect 42480 -27332 42538 -27074
rect 41174 -27334 42538 -27332
rect 41174 -27388 41186 -27334
rect 41962 -27388 42538 -27334
rect 41174 -27390 42538 -27388
rect 41174 -27395 41974 -27390
rect 41174 -27490 41974 -27485
rect 39978 -27492 41974 -27490
rect 39978 -27546 41186 -27492
rect 41962 -27546 41974 -27492
rect 39978 -27548 41974 -27546
rect 39978 -27806 40578 -27548
rect 41174 -27553 41974 -27548
rect 41174 -27648 41974 -27643
rect 42480 -27648 42538 -27390
rect 41174 -27650 42538 -27648
rect 41174 -27704 41186 -27650
rect 41962 -27704 42538 -27650
rect 41174 -27706 42538 -27704
rect 41174 -27711 41974 -27706
rect 41174 -27806 41974 -27801
rect 39978 -27808 41974 -27806
rect 39978 -27862 41186 -27808
rect 41962 -27862 41974 -27808
rect 39978 -27864 41974 -27862
rect 39978 -28122 40578 -27864
rect 41174 -27869 41974 -27864
rect 41174 -27964 41974 -27959
rect 42480 -27964 42538 -27706
rect 41174 -27966 42538 -27964
rect 41174 -28020 41186 -27966
rect 41962 -28020 42538 -27966
rect 41174 -28022 42538 -28020
rect 41174 -28027 41974 -28022
rect 41174 -28122 41974 -28117
rect 39978 -28124 41974 -28122
rect 39978 -28178 41186 -28124
rect 41962 -28178 41974 -28124
rect 39978 -28180 41974 -28178
rect 39978 -28438 40578 -28180
rect 41174 -28185 41974 -28180
rect 41174 -28280 41974 -28275
rect 42480 -28280 42538 -28022
rect 41174 -28282 42538 -28280
rect 41174 -28336 41186 -28282
rect 41962 -28336 42538 -28282
rect 41174 -28338 42538 -28336
rect 41174 -28343 41974 -28338
rect 41174 -28438 41974 -28433
rect 39978 -28440 41974 -28438
rect 39978 -28494 41186 -28440
rect 41962 -28494 41974 -28440
rect 39978 -28496 41974 -28494
rect 39978 -28754 40578 -28496
rect 41174 -28501 41974 -28496
rect 41174 -28596 41974 -28591
rect 42480 -28596 42538 -28338
rect 41174 -28598 42538 -28596
rect 41174 -28652 41186 -28598
rect 41962 -28652 42538 -28598
rect 41174 -28654 42538 -28652
rect 41174 -28659 41974 -28654
rect 41174 -28754 41974 -28749
rect 39978 -28756 41974 -28754
rect 39978 -28810 41186 -28756
rect 41962 -28810 41974 -28756
rect 39978 -28812 41974 -28810
rect 39978 -29070 40578 -28812
rect 41174 -28817 41974 -28812
rect 41174 -28912 41974 -28907
rect 42480 -28912 42538 -28654
rect 41174 -28914 42538 -28912
rect 41174 -28968 41186 -28914
rect 41962 -28968 42538 -28914
rect 41174 -28970 42538 -28968
rect 41174 -28975 41974 -28970
rect 41174 -29070 41974 -29065
rect 39978 -29072 41974 -29070
rect 39978 -29126 41186 -29072
rect 41962 -29126 41974 -29072
rect 39978 -29128 41974 -29126
rect 39978 -29386 40578 -29128
rect 41174 -29133 41974 -29128
rect 41174 -29228 41974 -29223
rect 42480 -29228 42538 -28970
rect 41174 -29230 42538 -29228
rect 41174 -29284 41186 -29230
rect 41962 -29284 42538 -29230
rect 41174 -29286 42538 -29284
rect 41174 -29291 41974 -29286
rect 41174 -29386 41974 -29381
rect 39978 -29388 41974 -29386
rect 39978 -29442 41186 -29388
rect 41962 -29442 41974 -29388
rect 39978 -29444 41974 -29442
rect 39978 -29702 40578 -29444
rect 41174 -29449 41974 -29444
rect 41174 -29544 41974 -29539
rect 42480 -29544 42538 -29286
rect 41174 -29546 42538 -29544
rect 41174 -29600 41186 -29546
rect 41962 -29600 42538 -29546
rect 41174 -29602 42538 -29600
rect 41174 -29607 41974 -29602
rect 41174 -29702 41974 -29697
rect 39978 -29704 41974 -29702
rect 39978 -29758 41186 -29704
rect 41962 -29758 41974 -29704
rect 39978 -29760 41974 -29758
rect 39978 -30018 40578 -29760
rect 41174 -29765 41974 -29760
rect 41174 -29860 41974 -29855
rect 42480 -29860 42538 -29602
rect 41174 -29862 42538 -29860
rect 41174 -29916 41186 -29862
rect 41962 -29916 42538 -29862
rect 41174 -29918 42538 -29916
rect 41174 -29923 41974 -29918
rect 41174 -30018 41974 -30013
rect 39978 -30020 41974 -30018
rect 39978 -30074 41186 -30020
rect 41962 -30074 41974 -30020
rect 39978 -30076 41974 -30074
rect 39978 -30334 40578 -30076
rect 41174 -30081 41974 -30076
rect 41174 -30176 41974 -30171
rect 42480 -30176 42538 -29918
rect 41174 -30178 42538 -30176
rect 41174 -30232 41186 -30178
rect 41962 -30232 42538 -30178
rect 41174 -30234 42538 -30232
rect 41174 -30239 41974 -30234
rect 41174 -30334 41974 -30329
rect 39978 -30336 41974 -30334
rect 39978 -30390 41186 -30336
rect 41962 -30390 41974 -30336
rect 39978 -30392 41974 -30390
rect 3976 -30482 4399 -30470
rect -4155 -30876 -3272 -30759
rect -4155 -30878 -3941 -30876
rect -4397 -31444 -3941 -30878
rect -3373 -30878 -1892 -30876
rect -3373 -31444 1204 -30878
rect 3976 -30882 3988 -30482
rect 4388 -30882 4399 -30482
rect 3976 -30893 4399 -30882
rect 39978 -30650 40578 -30392
rect 41174 -30397 41974 -30392
rect 41174 -30492 41974 -30487
rect 42480 -30492 42538 -30234
rect 41174 -30494 42538 -30492
rect 41174 -30548 41186 -30494
rect 41962 -30548 42538 -30494
rect 41174 -30550 42538 -30548
rect 41174 -30555 41974 -30550
rect 41174 -30650 41974 -30645
rect 39978 -30652 41974 -30650
rect 39978 -30706 41186 -30652
rect 41962 -30706 41974 -30652
rect 39978 -30708 41974 -30706
rect -4155 -31608 -3272 -31444
rect 636 -31523 1204 -31444
rect 636 -31621 3374 -31523
rect 636 -31656 1974 -31621
rect 636 -31729 642 -31656
rect 1967 -31729 1974 -31656
rect 636 -31735 1974 -31729
rect 636 -31875 694 -31735
rect 636 -32862 639 -31875
rect 692 -32862 694 -31875
rect 636 -32868 694 -32862
rect 764 -31875 822 -31868
rect 764 -32862 767 -31875
rect 820 -32862 822 -31875
rect 360 -32903 432 -32898
rect 360 -32909 682 -32903
rect 360 -32912 620 -32909
rect 360 -32968 368 -32912
rect 424 -32965 620 -32912
rect 676 -32965 682 -32909
rect 424 -32968 682 -32965
rect 360 -32971 682 -32968
rect 360 -32974 432 -32971
rect -1245 -33020 -785 -32990
rect 764 -33020 822 -32862
rect 892 -31875 950 -31735
rect 892 -32862 895 -31875
rect 948 -32862 950 -31875
rect 892 -32868 950 -32862
rect 1020 -31875 1078 -31868
rect 1020 -32862 1023 -31875
rect 1076 -32862 1078 -31875
rect 1020 -33020 1078 -32862
rect 1148 -31875 1206 -31735
rect 1148 -32862 1151 -31875
rect 1204 -32862 1206 -31875
rect 1148 -32868 1206 -32862
rect 1276 -31875 1334 -31868
rect 1276 -32862 1279 -31875
rect 1332 -32862 1334 -31875
rect 1276 -33020 1334 -32862
rect 1404 -31875 1462 -31735
rect 1404 -32862 1407 -31875
rect 1460 -32862 1462 -31875
rect 1404 -32868 1462 -32862
rect 1532 -31875 1590 -31868
rect 1532 -32862 1535 -31875
rect 1588 -32862 1590 -31875
rect 1532 -33020 1590 -32862
rect 1660 -31875 1718 -31735
rect 1660 -32862 1663 -31875
rect 1716 -32862 1718 -31875
rect 1660 -32868 1718 -32862
rect 1788 -31875 1846 -31868
rect 1788 -32862 1791 -31875
rect 1844 -32862 1846 -31875
rect 1788 -33020 1846 -32862
rect 1916 -31875 1974 -31735
rect 1916 -32862 1919 -31875
rect 1972 -32862 1974 -31875
rect 1916 -32868 1974 -32862
rect 2348 -32473 2414 -31621
rect 2540 -32473 2606 -31621
rect 2732 -32473 2798 -31621
rect 2924 -32473 2990 -31621
rect 3116 -32473 3182 -31621
rect 3308 -32473 3374 -31621
rect 3541 -31888 3646 -31863
rect 3541 -31944 3563 -31888
rect 3619 -31944 3646 -31888
rect 3541 -31961 3646 -31944
rect 2348 -32867 2354 -32473
rect 2408 -32867 2414 -32473
rect 2348 -32873 2414 -32867
rect 2444 -32867 2450 -32473
rect 2504 -32867 2510 -32473
rect 1904 -32907 2396 -32901
rect 1904 -32909 1911 -32907
rect 1896 -32960 1911 -32909
rect 1983 -32908 2396 -32907
rect 1983 -32960 2338 -32908
rect 1896 -32961 2338 -32960
rect 2390 -32961 2396 -32908
rect 1896 -32965 2396 -32961
rect 2332 -32967 2396 -32965
rect 2444 -33011 2510 -32867
rect 2540 -32867 2546 -32473
rect 2600 -32867 2606 -32473
rect 2540 -32873 2606 -32867
rect 2636 -32867 2642 -32473
rect 2696 -32867 2702 -32473
rect 2636 -33011 2702 -32867
rect 2732 -32867 2738 -32473
rect 2792 -32867 2798 -32473
rect 2732 -32873 2798 -32867
rect 2828 -32867 2834 -32473
rect 2888 -32867 2894 -32473
rect 2828 -33011 2894 -32867
rect 2924 -32867 2930 -32473
rect 2984 -32867 2990 -32473
rect 2924 -32873 2990 -32867
rect 3020 -32867 3026 -32473
rect 3080 -32867 3086 -32473
rect 3020 -33011 3086 -32867
rect 3116 -32867 3122 -32473
rect 3176 -32867 3182 -32473
rect 3116 -32873 3182 -32867
rect 3212 -32867 3218 -32473
rect 3272 -32867 3278 -32473
rect 3212 -33011 3278 -32867
rect 3308 -32867 3314 -32473
rect 3368 -32867 3374 -32473
rect 3308 -32873 3374 -32867
rect 3558 -32901 3628 -31961
rect 3314 -32907 3628 -32901
rect 3314 -32963 3320 -32907
rect 3390 -32963 3628 -32907
rect 3314 -32971 3628 -32963
rect 3988 -33011 4388 -30893
rect -1245 -33420 -1215 -33020
rect -815 -33420 1846 -33020
rect 2443 -33411 4388 -33011
rect 39978 -30966 40578 -30708
rect 41174 -30713 41974 -30708
rect 41174 -30808 41974 -30803
rect 42480 -30808 42538 -30550
rect 41174 -30810 42538 -30808
rect 41174 -30864 41186 -30810
rect 41962 -30864 42538 -30810
rect 41174 -30866 42538 -30864
rect 41174 -30871 41974 -30866
rect 41174 -30966 41974 -30961
rect 39978 -30968 41974 -30966
rect 39978 -31022 41186 -30968
rect 41962 -31022 41974 -30968
rect 39978 -31024 41974 -31022
rect 39978 -31282 40578 -31024
rect 41174 -31029 41974 -31024
rect 41174 -31124 41974 -31119
rect 42480 -31124 42538 -30866
rect 41174 -31126 42538 -31124
rect 41174 -31180 41186 -31126
rect 41962 -31180 42538 -31126
rect 41174 -31182 42538 -31180
rect 41174 -31187 41974 -31182
rect 41174 -31282 41974 -31277
rect 39978 -31284 41974 -31282
rect 39978 -31338 41186 -31284
rect 41962 -31338 41974 -31284
rect 39978 -31340 41974 -31338
rect 39978 -31598 40578 -31340
rect 41174 -31345 41974 -31340
rect 41174 -31440 41974 -31435
rect 42480 -31440 42538 -31182
rect 41174 -31442 42538 -31440
rect 41174 -31496 41186 -31442
rect 41962 -31496 42538 -31442
rect 41174 -31498 42538 -31496
rect 41174 -31503 41974 -31498
rect 41174 -31598 41974 -31593
rect 39978 -31600 41974 -31598
rect 39978 -31654 41186 -31600
rect 41962 -31654 41974 -31600
rect 39978 -31656 41974 -31654
rect 39978 -31914 40578 -31656
rect 41174 -31661 41974 -31656
rect 41174 -31756 41974 -31751
rect 42480 -31756 42538 -31498
rect 41174 -31758 42538 -31756
rect 41174 -31812 41186 -31758
rect 41962 -31812 42538 -31758
rect 41174 -31814 42538 -31812
rect 41174 -31819 41974 -31814
rect 41174 -31914 41974 -31909
rect 39978 -31916 41974 -31914
rect 39978 -31970 41186 -31916
rect 41962 -31970 41974 -31916
rect 39978 -31972 41974 -31970
rect 39978 -32230 40578 -31972
rect 41174 -31977 41974 -31972
rect 41174 -32072 41974 -32067
rect 42480 -32072 42538 -31814
rect 41174 -32074 42538 -32072
rect 41174 -32128 41186 -32074
rect 41962 -32128 42538 -32074
rect 41174 -32130 42538 -32128
rect 41174 -32135 41974 -32130
rect 41174 -32230 41974 -32225
rect 39978 -32232 41974 -32230
rect 39978 -32286 41186 -32232
rect 41962 -32286 41974 -32232
rect 39978 -32288 41974 -32286
rect 39978 -32546 40578 -32288
rect 41174 -32293 41974 -32288
rect 41174 -32388 41974 -32383
rect 42480 -32388 42538 -32130
rect 41174 -32390 42538 -32388
rect 41174 -32444 41186 -32390
rect 41962 -32444 42538 -32390
rect 41174 -32446 42538 -32444
rect 41174 -32451 41974 -32446
rect 41174 -32546 41974 -32541
rect 39978 -32548 41974 -32546
rect 39978 -32602 41186 -32548
rect 41962 -32602 41974 -32548
rect 39978 -32604 41974 -32602
rect 39978 -32862 40578 -32604
rect 41174 -32609 41974 -32604
rect 41174 -32704 41974 -32699
rect 42480 -32704 42538 -32446
rect 41174 -32706 42538 -32704
rect 41174 -32760 41186 -32706
rect 41962 -32760 42538 -32706
rect 41174 -32762 42538 -32760
rect 41174 -32767 41974 -32762
rect 41174 -32862 41974 -32857
rect 39978 -32864 41974 -32862
rect 39978 -32918 41186 -32864
rect 41962 -32918 41974 -32864
rect 39978 -32920 41974 -32918
rect 39978 -33178 40578 -32920
rect 41174 -32925 41974 -32920
rect 41174 -33020 41974 -33015
rect 42480 -33020 42538 -32762
rect 41174 -33022 42538 -33020
rect 41174 -33076 41186 -33022
rect 41962 -33076 42538 -33022
rect 41174 -33078 42538 -33076
rect 41174 -33083 41974 -33078
rect 41174 -33178 41974 -33173
rect 39978 -33180 41974 -33178
rect 39978 -33234 41186 -33180
rect 41962 -33234 41974 -33180
rect 39978 -33236 41974 -33234
rect -1245 -33450 -785 -33420
rect 636 -33567 694 -33560
rect 636 -34554 639 -33567
rect 692 -34554 694 -33567
rect 636 -34809 694 -34554
rect 764 -33567 822 -33420
rect 764 -34554 767 -33567
rect 820 -34554 822 -33567
rect 764 -34560 822 -34554
rect 892 -33567 950 -33560
rect 892 -34554 895 -33567
rect 948 -34554 950 -33567
rect 892 -34809 950 -34554
rect 1020 -33567 1078 -33420
rect 1020 -34554 1023 -33567
rect 1076 -34554 1078 -33567
rect 1020 -34560 1078 -34554
rect 1148 -33567 1206 -33560
rect 1148 -34554 1151 -33567
rect 1204 -34554 1206 -33567
rect 1148 -34809 1206 -34554
rect 1276 -33567 1334 -33420
rect 1276 -34554 1279 -33567
rect 1332 -34554 1334 -33567
rect 1276 -34560 1334 -34554
rect 1404 -33567 1462 -33560
rect 1404 -34554 1407 -33567
rect 1460 -34554 1462 -33567
rect 1404 -34809 1462 -34554
rect 1532 -33567 1590 -33420
rect 1532 -34554 1535 -33567
rect 1588 -34554 1590 -33567
rect 1532 -34560 1590 -34554
rect 1660 -33567 1718 -33560
rect 1660 -34554 1663 -33567
rect 1716 -34554 1718 -33567
rect 1660 -34809 1718 -34554
rect 1788 -33567 1846 -33420
rect 2324 -33455 2409 -33454
rect 1902 -33460 2409 -33455
rect 1902 -33461 2331 -33460
rect 1902 -33514 1909 -33461
rect 1981 -33513 2331 -33461
rect 2403 -33513 2409 -33460
rect 1981 -33514 2409 -33513
rect 1902 -33519 2409 -33514
rect 1788 -34554 1791 -33567
rect 1844 -34554 1846 -33567
rect 1788 -34560 1846 -34554
rect 1916 -33567 1974 -33560
rect 1916 -34554 1919 -33567
rect 1972 -34554 1974 -33567
rect 2444 -34351 2508 -33411
rect 2636 -34351 2700 -33411
rect 2828 -34351 2892 -33411
rect 3020 -34351 3084 -33411
rect 3212 -34351 3276 -33411
rect 39978 -33494 40578 -33236
rect 41174 -33241 41974 -33236
rect 41174 -33336 41974 -33331
rect 42480 -33336 42538 -33078
rect 41174 -33338 42538 -33336
rect 41174 -33392 41186 -33338
rect 41962 -33392 42538 -33338
rect 41174 -33394 42538 -33392
rect 41174 -33399 41974 -33394
rect 41174 -33494 41974 -33489
rect 39978 -33496 41974 -33494
rect 39978 -33550 41186 -33496
rect 41962 -33550 41974 -33496
rect 39978 -33552 41974 -33550
rect 3312 -33770 3838 -33757
rect 3312 -33776 3683 -33770
rect 3312 -33909 3322 -33776
rect 3374 -33909 3683 -33776
rect 3822 -33909 3838 -33770
rect 3312 -33923 3838 -33909
rect 39978 -33810 40578 -33552
rect 41174 -33557 41974 -33552
rect 41174 -33652 41974 -33647
rect 42480 -33652 42538 -33394
rect 41174 -33654 42538 -33652
rect 41174 -33708 41186 -33654
rect 41962 -33708 42538 -33654
rect 41174 -33710 42538 -33708
rect 41174 -33715 41974 -33710
rect 41174 -33810 41974 -33805
rect 39978 -33812 41974 -33810
rect 39978 -33866 41186 -33812
rect 41962 -33866 41974 -33812
rect 39978 -33868 41974 -33866
rect 39978 -34126 40578 -33868
rect 41174 -33873 41974 -33868
rect 41174 -33968 41974 -33963
rect 42480 -33968 42538 -33710
rect 41174 -33970 42538 -33968
rect 41174 -34024 41186 -33970
rect 41962 -34024 42538 -33970
rect 41174 -34026 42538 -34024
rect 41174 -34031 41974 -34026
rect 41174 -34126 41974 -34121
rect 39978 -34128 41974 -34126
rect 39978 -34182 41186 -34128
rect 41962 -34182 41974 -34128
rect 39978 -34184 41974 -34182
rect 1916 -34809 1974 -34554
rect -6172 -35150 -5411 -34864
rect -6172 -35536 -6013 -35150
rect -5627 -35536 -5411 -35150
rect -6172 -35739 -5411 -35536
rect 636 -35331 1974 -34809
rect 2348 -34545 2354 -34351
rect 2408 -34545 2414 -34351
rect 2348 -34671 2414 -34545
rect 2444 -34545 2450 -34351
rect 2504 -34545 2510 -34351
rect 2444 -34551 2510 -34545
rect 2540 -34545 2546 -34351
rect 2600 -34545 2606 -34351
rect 2540 -34671 2606 -34545
rect 2636 -34545 2642 -34351
rect 2696 -34545 2702 -34351
rect 2636 -34551 2702 -34545
rect 2732 -34545 2738 -34351
rect 2792 -34545 2798 -34351
rect 2732 -34671 2798 -34545
rect 2828 -34545 2834 -34351
rect 2888 -34545 2894 -34351
rect 2828 -34551 2894 -34545
rect 2924 -34545 2930 -34351
rect 2984 -34545 2990 -34351
rect 2924 -34671 2990 -34545
rect 3020 -34545 3026 -34351
rect 3080 -34545 3086 -34351
rect 3020 -34551 3086 -34545
rect 3116 -34545 3122 -34351
rect 3176 -34545 3182 -34351
rect 3116 -34671 3182 -34545
rect 3212 -34545 3218 -34351
rect 3272 -34545 3278 -34351
rect 3212 -34551 3278 -34545
rect 3308 -34545 3314 -34351
rect 3368 -34545 3374 -34351
rect 3308 -34671 3374 -34545
rect 2348 -34677 3374 -34671
rect 2348 -34755 2354 -34677
rect 2792 -34755 2930 -34677
rect 3368 -34755 3374 -34677
rect 2348 -34988 3374 -34755
rect 2348 -35150 2391 -34988
rect 3339 -35150 3374 -34988
rect 2348 -35176 3374 -35150
rect 39978 -34442 40578 -34184
rect 41174 -34189 41974 -34184
rect 41174 -34284 41974 -34279
rect 42480 -34284 42538 -34026
rect 41174 -34286 42538 -34284
rect 41174 -34340 41186 -34286
rect 41962 -34340 42538 -34286
rect 41174 -34342 42538 -34340
rect 41174 -34347 41974 -34342
rect 41174 -34442 41974 -34437
rect 39978 -34444 41974 -34442
rect 39978 -34498 41186 -34444
rect 41962 -34498 41974 -34444
rect 39978 -34500 41974 -34498
rect 39978 -34758 40578 -34500
rect 41174 -34505 41974 -34500
rect 41174 -34600 41974 -34595
rect 42480 -34600 42538 -34342
rect 41174 -34602 42538 -34600
rect 41174 -34656 41186 -34602
rect 41962 -34656 42538 -34602
rect 41174 -34658 42538 -34656
rect 41174 -34663 41974 -34658
rect 41174 -34758 41974 -34753
rect 39978 -34760 41974 -34758
rect 39978 -34814 41186 -34760
rect 41962 -34814 41974 -34760
rect 39978 -34816 41974 -34814
rect 39978 -35074 40578 -34816
rect 41174 -34821 41974 -34816
rect 41174 -34916 41974 -34911
rect 42480 -34916 42538 -34658
rect 41174 -34918 42538 -34916
rect 41174 -34972 41186 -34918
rect 41962 -34972 42538 -34918
rect 41174 -34974 42538 -34972
rect 41174 -34979 41974 -34974
rect 41174 -35074 41974 -35069
rect 39978 -35076 41974 -35074
rect 39978 -35130 41186 -35076
rect 41962 -35130 41974 -35076
rect 39978 -35132 41974 -35130
rect 39978 -35331 40578 -35132
rect 41174 -35137 41974 -35132
rect 41174 -35232 41974 -35227
rect 42480 -35232 42538 -34974
rect 41174 -35234 42538 -35232
rect 41174 -35288 41186 -35234
rect 41962 -35288 42538 -35234
rect 41174 -35290 42538 -35288
rect 41174 -35295 41974 -35290
rect 636 -35390 40578 -35331
rect 41174 -35390 41974 -35385
rect 636 -35392 41974 -35390
rect 636 -35446 41186 -35392
rect 41962 -35446 41974 -35392
rect 636 -35448 41974 -35446
rect 636 -35706 40578 -35448
rect 41174 -35453 41974 -35448
rect 41174 -35548 41974 -35543
rect 42480 -35548 42538 -35290
rect 41174 -35550 42538 -35548
rect 41174 -35604 41186 -35550
rect 41962 -35604 42538 -35550
rect 41174 -35606 42538 -35604
rect 41174 -35611 41974 -35606
rect 41174 -35706 41974 -35701
rect 636 -35708 41974 -35706
rect 636 -35762 41186 -35708
rect 41962 -35762 41974 -35708
rect 636 -35764 41974 -35762
rect 636 -35931 40578 -35764
rect 41174 -35769 41974 -35764
rect 41174 -35864 41974 -35859
rect 42480 -35864 42538 -35606
rect 41174 -35866 42538 -35864
rect 41174 -35920 41186 -35866
rect 41962 -35920 42538 -35866
rect 41174 -35922 42538 -35920
rect 41174 -35927 41974 -35922
rect 39978 -36022 40578 -35931
rect 41174 -36022 41974 -36017
rect 39978 -36024 41974 -36022
rect 39978 -36078 41186 -36024
rect 41962 -36078 41974 -36024
rect 39978 -36080 41974 -36078
rect 39978 -36338 40578 -36080
rect 41174 -36085 41974 -36080
rect 41174 -36180 41974 -36175
rect 42480 -36180 42538 -35922
rect 41174 -36182 42538 -36180
rect 41174 -36236 41186 -36182
rect 41962 -36236 42538 -36182
rect 41174 -36238 42538 -36236
rect 41174 -36243 41974 -36238
rect 41174 -36338 41974 -36333
rect 39978 -36340 41974 -36338
rect 39978 -36394 41186 -36340
rect 41962 -36394 41974 -36340
rect 39978 -36396 41974 -36394
rect 39978 -36654 40578 -36396
rect 41174 -36401 41974 -36396
rect 41174 -36496 41974 -36491
rect 42480 -36496 42538 -36238
rect 41174 -36498 42538 -36496
rect 41174 -36552 41186 -36498
rect 41962 -36552 42538 -36498
rect 41174 -36554 42538 -36552
rect 41174 -36559 41974 -36554
rect 41174 -36654 41974 -36649
rect 39978 -36656 41974 -36654
rect 39978 -36710 41186 -36656
rect 41962 -36710 41974 -36656
rect 39978 -36712 41974 -36710
rect 39978 -36970 40578 -36712
rect 41174 -36717 41974 -36712
rect 41174 -36812 41974 -36807
rect 42480 -36812 42538 -36554
rect 41174 -36814 42538 -36812
rect 41174 -36868 41186 -36814
rect 41962 -36868 42538 -36814
rect 41174 -36870 42538 -36868
rect 41174 -36875 41974 -36870
rect 41174 -36970 41974 -36965
rect 39978 -36972 41974 -36970
rect 39978 -37026 41186 -36972
rect 41962 -37026 41974 -36972
rect 39978 -37028 41974 -37026
rect 39978 -37286 40578 -37028
rect 41174 -37033 41974 -37028
rect 41174 -37128 41974 -37123
rect 42480 -37128 42538 -36870
rect 41174 -37130 42538 -37128
rect 41174 -37184 41186 -37130
rect 41962 -37184 42538 -37130
rect 41174 -37186 42538 -37184
rect 41174 -37191 41974 -37186
rect 41174 -37286 41974 -37281
rect 39978 -37288 41974 -37286
rect 39978 -37342 41186 -37288
rect 41962 -37342 41974 -37288
rect 39978 -37344 41974 -37342
rect 39978 -37602 40578 -37344
rect 41174 -37349 41974 -37344
rect 41174 -37444 41974 -37439
rect 42480 -37444 42538 -37186
rect 41174 -37446 42538 -37444
rect 41174 -37500 41186 -37446
rect 41962 -37500 42538 -37446
rect 41174 -37502 42538 -37500
rect 41174 -37507 41974 -37502
rect 41174 -37602 41974 -37597
rect 39978 -37604 41974 -37602
rect 39978 -37658 41186 -37604
rect 41962 -37658 41974 -37604
rect 39978 -37660 41974 -37658
rect 39978 -37918 40578 -37660
rect 41174 -37665 41974 -37660
rect 41174 -37760 41974 -37755
rect 42480 -37760 42538 -37502
rect 41174 -37762 42538 -37760
rect 41174 -37816 41186 -37762
rect 41962 -37816 42538 -37762
rect 41174 -37818 42538 -37816
rect 41174 -37823 41974 -37818
rect 41174 -37918 41974 -37913
rect 39978 -37920 41974 -37918
rect 39978 -37974 41186 -37920
rect 41962 -37974 41974 -37920
rect 39978 -37976 41974 -37974
rect 39978 -38234 40578 -37976
rect 41174 -37981 41974 -37976
rect 41174 -38076 41974 -38071
rect 42480 -38076 42538 -37818
rect 41174 -38078 42538 -38076
rect 41174 -38132 41186 -38078
rect 41962 -38132 42538 -38078
rect 41174 -38134 42538 -38132
rect 41174 -38139 41974 -38134
rect 41174 -38234 41974 -38229
rect 39978 -38236 41974 -38234
rect 39978 -38290 41186 -38236
rect 41962 -38290 41974 -38236
rect 39978 -38292 41974 -38290
rect 39978 -38550 40578 -38292
rect 41174 -38297 41974 -38292
rect 41174 -38392 41974 -38387
rect 42480 -38392 42538 -38134
rect 41174 -38394 42538 -38392
rect 41174 -38448 41186 -38394
rect 41962 -38448 42538 -38394
rect 41174 -38450 42538 -38448
rect 41174 -38455 41974 -38450
rect 41174 -38550 41974 -38545
rect 39978 -38552 41974 -38550
rect 39978 -38606 41186 -38552
rect 41962 -38606 41974 -38552
rect 39978 -38608 41974 -38606
rect 3976 -44482 4399 -44470
rect -4155 -44876 -3272 -44759
rect -4155 -45444 -3941 -44876
rect -3373 -44878 -1892 -44876
rect -3373 -45444 1204 -44878
rect 3976 -44882 3988 -44482
rect 4388 -44882 4399 -44482
rect 3976 -44893 4399 -44882
rect -4155 -45608 -3272 -45444
rect 636 -45523 1204 -45444
rect 636 -45621 3374 -45523
rect 636 -45656 1974 -45621
rect 636 -45729 642 -45656
rect 1967 -45729 1974 -45656
rect 636 -45735 1974 -45729
rect 636 -45875 694 -45735
rect 636 -46862 639 -45875
rect 692 -46862 694 -45875
rect 636 -46868 694 -46862
rect 764 -45875 822 -45868
rect 764 -46862 767 -45875
rect 820 -46862 822 -45875
rect 360 -46903 432 -46898
rect 360 -46909 682 -46903
rect 360 -46912 620 -46909
rect 360 -46968 368 -46912
rect 424 -46965 620 -46912
rect 676 -46965 682 -46909
rect 424 -46968 682 -46965
rect 360 -46971 682 -46968
rect 360 -46974 432 -46971
rect -1245 -47020 -785 -46990
rect 764 -47020 822 -46862
rect 892 -45875 950 -45735
rect 892 -46862 895 -45875
rect 948 -46862 950 -45875
rect 892 -46868 950 -46862
rect 1020 -45875 1078 -45868
rect 1020 -46862 1023 -45875
rect 1076 -46862 1078 -45875
rect 1020 -47020 1078 -46862
rect 1148 -45875 1206 -45735
rect 1148 -46862 1151 -45875
rect 1204 -46862 1206 -45875
rect 1148 -46868 1206 -46862
rect 1276 -45875 1334 -45868
rect 1276 -46862 1279 -45875
rect 1332 -46862 1334 -45875
rect 1276 -47020 1334 -46862
rect 1404 -45875 1462 -45735
rect 1404 -46862 1407 -45875
rect 1460 -46862 1462 -45875
rect 1404 -46868 1462 -46862
rect 1532 -45875 1590 -45868
rect 1532 -46862 1535 -45875
rect 1588 -46862 1590 -45875
rect 1532 -47020 1590 -46862
rect 1660 -45875 1718 -45735
rect 1660 -46862 1663 -45875
rect 1716 -46862 1718 -45875
rect 1660 -46868 1718 -46862
rect 1788 -45875 1846 -45868
rect 1788 -46862 1791 -45875
rect 1844 -46862 1846 -45875
rect 1788 -47020 1846 -46862
rect 1916 -45875 1974 -45735
rect 1916 -46862 1919 -45875
rect 1972 -46862 1974 -45875
rect 1916 -46868 1974 -46862
rect 2348 -46473 2414 -45621
rect 2540 -46473 2606 -45621
rect 2732 -46473 2798 -45621
rect 2924 -46473 2990 -45621
rect 3116 -46473 3182 -45621
rect 3308 -46473 3374 -45621
rect 3541 -45888 3646 -45863
rect 3541 -45944 3563 -45888
rect 3619 -45944 3646 -45888
rect 3541 -45961 3646 -45944
rect 2348 -46867 2354 -46473
rect 2408 -46867 2414 -46473
rect 2348 -46873 2414 -46867
rect 2444 -46867 2450 -46473
rect 2504 -46867 2510 -46473
rect 1904 -46907 2396 -46901
rect 1904 -46909 1911 -46907
rect 1896 -46960 1911 -46909
rect 1983 -46908 2396 -46907
rect 1983 -46960 2338 -46908
rect 1896 -46961 2338 -46960
rect 2390 -46961 2396 -46908
rect 1896 -46965 2396 -46961
rect 2332 -46967 2396 -46965
rect 2444 -47011 2510 -46867
rect 2540 -46867 2546 -46473
rect 2600 -46867 2606 -46473
rect 2540 -46873 2606 -46867
rect 2636 -46867 2642 -46473
rect 2696 -46867 2702 -46473
rect 2636 -47011 2702 -46867
rect 2732 -46867 2738 -46473
rect 2792 -46867 2798 -46473
rect 2732 -46873 2798 -46867
rect 2828 -46867 2834 -46473
rect 2888 -46867 2894 -46473
rect 2828 -47011 2894 -46867
rect 2924 -46867 2930 -46473
rect 2984 -46867 2990 -46473
rect 2924 -46873 2990 -46867
rect 3020 -46867 3026 -46473
rect 3080 -46867 3086 -46473
rect 3020 -47011 3086 -46867
rect 3116 -46867 3122 -46473
rect 3176 -46867 3182 -46473
rect 3116 -46873 3182 -46867
rect 3212 -46867 3218 -46473
rect 3272 -46867 3278 -46473
rect 3212 -47011 3278 -46867
rect 3308 -46867 3314 -46473
rect 3368 -46867 3374 -46473
rect 3308 -46873 3374 -46867
rect 3558 -46901 3628 -45961
rect 3314 -46907 3628 -46901
rect 3314 -46963 3320 -46907
rect 3390 -46963 3628 -46907
rect 3314 -46971 3628 -46963
rect 3988 -47011 4388 -44893
rect -1245 -47420 -1215 -47020
rect -815 -47420 1846 -47020
rect 2443 -47411 4388 -47011
rect -1245 -47450 -785 -47420
rect 636 -47567 694 -47560
rect 636 -48554 639 -47567
rect 692 -48554 694 -47567
rect 636 -48809 694 -48554
rect 764 -47567 822 -47420
rect 764 -48554 767 -47567
rect 820 -48554 822 -47567
rect 764 -48560 822 -48554
rect 892 -47567 950 -47560
rect 892 -48554 895 -47567
rect 948 -48554 950 -47567
rect 892 -48809 950 -48554
rect 1020 -47567 1078 -47420
rect 1020 -48554 1023 -47567
rect 1076 -48554 1078 -47567
rect 1020 -48560 1078 -48554
rect 1148 -47567 1206 -47560
rect 1148 -48554 1151 -47567
rect 1204 -48554 1206 -47567
rect 1148 -48809 1206 -48554
rect 1276 -47567 1334 -47420
rect 1276 -48554 1279 -47567
rect 1332 -48554 1334 -47567
rect 1276 -48560 1334 -48554
rect 1404 -47567 1462 -47560
rect 1404 -48554 1407 -47567
rect 1460 -48554 1462 -47567
rect 1404 -48809 1462 -48554
rect 1532 -47567 1590 -47420
rect 1532 -48554 1535 -47567
rect 1588 -48554 1590 -47567
rect 1532 -48560 1590 -48554
rect 1660 -47567 1718 -47560
rect 1660 -48554 1663 -47567
rect 1716 -48554 1718 -47567
rect 1660 -48809 1718 -48554
rect 1788 -47567 1846 -47420
rect 2324 -47455 2409 -47454
rect 1902 -47460 2409 -47455
rect 1902 -47461 2331 -47460
rect 1902 -47514 1909 -47461
rect 1981 -47513 2331 -47461
rect 2403 -47513 2409 -47460
rect 1981 -47514 2409 -47513
rect 1902 -47519 2409 -47514
rect 1788 -48554 1791 -47567
rect 1844 -48554 1846 -47567
rect 1788 -48560 1846 -48554
rect 1916 -47567 1974 -47560
rect 1916 -48554 1919 -47567
rect 1972 -48554 1974 -47567
rect 2444 -48351 2508 -47411
rect 2636 -48351 2700 -47411
rect 2828 -48351 2892 -47411
rect 3020 -48351 3084 -47411
rect 3212 -48351 3276 -47411
rect 3312 -47770 3838 -47757
rect 3312 -47776 3683 -47770
rect 3312 -47909 3322 -47776
rect 3374 -47909 3683 -47776
rect 3822 -47909 3838 -47770
rect 3312 -47923 3838 -47909
rect 1916 -48809 1974 -48554
rect -6172 -49150 -5411 -48864
rect -6172 -49536 -6013 -49150
rect -5627 -49536 -5411 -49150
rect -6172 -49739 -5411 -49536
rect 636 -49331 1974 -48809
rect 2348 -48545 2354 -48351
rect 2408 -48545 2414 -48351
rect 2348 -48671 2414 -48545
rect 2444 -48545 2450 -48351
rect 2504 -48545 2510 -48351
rect 2444 -48551 2510 -48545
rect 2540 -48545 2546 -48351
rect 2600 -48545 2606 -48351
rect 2540 -48671 2606 -48545
rect 2636 -48545 2642 -48351
rect 2696 -48545 2702 -48351
rect 2636 -48551 2702 -48545
rect 2732 -48545 2738 -48351
rect 2792 -48545 2798 -48351
rect 2732 -48671 2798 -48545
rect 2828 -48545 2834 -48351
rect 2888 -48545 2894 -48351
rect 2828 -48551 2894 -48545
rect 2924 -48545 2930 -48351
rect 2984 -48545 2990 -48351
rect 2924 -48671 2990 -48545
rect 3020 -48545 3026 -48351
rect 3080 -48545 3086 -48351
rect 3020 -48551 3086 -48545
rect 3116 -48545 3122 -48351
rect 3176 -48545 3182 -48351
rect 3116 -48671 3182 -48545
rect 3212 -48545 3218 -48351
rect 3272 -48545 3278 -48351
rect 3212 -48551 3278 -48545
rect 3308 -48545 3314 -48351
rect 3368 -48545 3374 -48351
rect 3308 -48671 3374 -48545
rect 2348 -48677 3374 -48671
rect 2348 -48755 2354 -48677
rect 2792 -48755 2930 -48677
rect 3368 -48755 3374 -48677
rect 2348 -48988 3374 -48755
rect 2348 -49150 2391 -48988
rect 3339 -49150 3374 -48988
rect 2348 -49176 3374 -49150
rect 39978 -49331 40578 -38608
rect 41174 -38613 41974 -38608
rect 636 -49931 40578 -49331
<< via2 >>
rect -4014 1487 -3442 2059
rect -5966 -552 -5627 -213
rect 1065 -217 1136 -146
rect 879 -374 947 -306
rect 3753 -217 3824 -146
rect 3567 -374 3635 -306
rect -3941 -3444 -3373 -2876
rect 3988 -2882 4388 -2482
rect 12686 739 12778 831
rect 6441 -217 6512 -146
rect 6255 -374 6323 -306
rect 9129 -217 9200 -146
rect 8943 -374 9011 -306
rect 19140 400 19460 720
rect 18147 -1198 18235 -1110
rect 14612 -2636 14682 -2566
rect -1215 -5420 -815 -5020
rect -6013 -7536 -5627 -7150
rect 42450 -12096 42510 -12036
rect -3941 -17444 -3373 -16876
rect 4080 -16882 4388 -16482
rect -1215 -19420 -815 -19020
rect -6013 -21536 -5627 -21150
rect 41132 -25633 41320 -25445
rect 41053 -26151 41128 -26056
rect -3941 -31444 -3373 -30876
rect 3988 -30882 4388 -30482
rect -1215 -33420 -815 -33020
rect -6013 -35536 -5627 -35150
rect -3941 -45444 -3373 -44876
rect 3988 -44882 4388 -44482
rect -1215 -47420 -815 -47020
rect -6013 -49536 -5627 -49150
<< metal3 >>
rect -4072 2064 -3400 2092
rect -4072 1482 -4019 2064
rect -3437 1482 -3400 2064
rect -4072 1429 -3400 1482
rect 12540 836 12928 983
rect 12540 734 12681 836
rect 12783 734 12928 836
rect 12540 586 12928 734
rect 19038 720 19500 784
rect 19038 400 19140 720
rect 19460 400 19500 720
rect 19038 337 19500 400
rect -6127 -208 -5411 -70
rect 1208 -137 1297 -136
rect -6127 -557 -5971 -208
rect -5622 -557 -5411 -208
rect 1056 -146 9209 -137
rect 1056 -217 1065 -146
rect 1136 -217 3753 -146
rect 3824 -217 6441 -146
rect 6512 -217 9129 -146
rect 9200 -217 9209 -146
rect 1056 -226 9209 -217
rect 864 -301 962 -291
rect 864 -379 874 -301
rect 952 -379 962 -301
rect 864 -389 962 -379
rect -6127 -683 -5411 -557
rect -2070 -1034 -1654 -946
rect -2070 -1282 -1998 -1034
rect -1750 -1113 -1654 -1034
rect 1208 -1113 1297 -226
rect 3552 -301 3650 -291
rect 3552 -379 3562 -301
rect 3640 -379 3650 -301
rect 3552 -389 3650 -379
rect 6240 -301 6338 -291
rect 6240 -379 6250 -301
rect 6328 -379 6338 -301
rect 6240 -389 6338 -379
rect 8928 -301 9026 -291
rect 8928 -379 8938 -301
rect 9016 -379 9026 -301
rect 8928 -389 9026 -379
rect -1750 -1202 1297 -1113
rect 17925 -1042 18390 -929
rect 17925 -1105 41325 -1042
rect -1750 -1282 -1654 -1202
rect -2070 -1372 -1654 -1282
rect 17925 -1203 18142 -1105
rect 18240 -1203 41325 -1105
rect 17925 -1240 41325 -1203
rect 17925 -1367 18390 -1240
rect 3976 -2477 4399 -2470
rect -4155 -2871 -3272 -2759
rect -4155 -3449 -3946 -2871
rect -3368 -3449 -3272 -2871
rect 3976 -2887 3983 -2477
rect 4393 -2887 4399 -2477
rect 14607 -2566 14687 -2561
rect 14607 -2636 14612 -2566
rect 14682 -2636 40398 -2566
rect 40468 -2636 40474 -2566
rect 14607 -2641 14687 -2636
rect 3976 -2893 4399 -2887
rect -4155 -3608 -3272 -3449
rect -1245 -5015 -245 -4990
rect -1245 -5425 -1220 -5015
rect -810 -5425 -245 -5015
rect -1245 -5450 -245 -5425
rect -6172 -7145 -5411 -6864
rect -6172 -7541 -6018 -7145
rect -5622 -7541 -5411 -7145
rect -6172 -7739 -5411 -7541
rect 3976 -16477 4399 -16470
rect -4155 -16871 -3272 -16759
rect -4155 -17449 -3946 -16871
rect -3368 -17449 -3272 -16871
rect 3976 -16887 3983 -16477
rect 4393 -16887 4399 -16477
rect 3976 -16893 4399 -16887
rect -4155 -17608 -3272 -17449
rect -1245 -19015 -245 -18990
rect -1245 -19425 -1220 -19015
rect -810 -19425 -245 -19015
rect -1245 -19450 -245 -19425
rect -6172 -21145 -5411 -20864
rect -6172 -21541 -6018 -21145
rect -5622 -21541 -5411 -21145
rect -6172 -21739 -5411 -21541
rect 41127 -25417 41325 -1240
rect 42425 -12032 42537 -12016
rect 42425 -12100 42446 -12032
rect 42514 -12100 42537 -12032
rect 42425 -12114 42537 -12100
rect 41007 -25445 41349 -25417
rect 41007 -25633 41132 -25445
rect 41320 -25633 41349 -25445
rect 41007 -25654 41349 -25633
rect 41007 -26056 41147 -25654
rect 41007 -26151 41053 -26056
rect 41128 -26151 41147 -26056
rect 41007 -26171 41147 -26151
rect 3976 -30477 4399 -30470
rect -4155 -30871 -3272 -30759
rect -4155 -31449 -3946 -30871
rect -3368 -31449 -3272 -30871
rect 3976 -30887 3983 -30477
rect 4393 -30887 4399 -30477
rect 3976 -30893 4399 -30887
rect -4155 -31608 -3272 -31449
rect -1245 -33015 -245 -32990
rect -1245 -33425 -1220 -33015
rect -810 -33425 -245 -33015
rect -1245 -33450 -245 -33425
rect -6172 -35145 -5411 -34864
rect -6172 -35541 -6018 -35145
rect -5622 -35541 -5411 -35145
rect -6172 -35739 -5411 -35541
rect 3976 -44477 4399 -44470
rect -4155 -44871 -3272 -44759
rect -4155 -45449 -3946 -44871
rect -3368 -45449 -3272 -44871
rect 3976 -44887 3983 -44477
rect 4393 -44887 4399 -44477
rect 3976 -44893 4399 -44887
rect -4155 -45608 -3272 -45449
rect -1245 -47015 -245 -46990
rect -1245 -47425 -1220 -47015
rect -810 -47425 -245 -47015
rect -1245 -47450 -245 -47425
rect -6172 -49145 -5411 -48864
rect -6172 -49541 -6018 -49145
rect -5622 -49541 -5411 -49145
rect -6172 -49739 -5411 -49541
<< via3 >>
rect -4019 2059 -3437 2064
rect -4019 1487 -4014 2059
rect -4014 1487 -3442 2059
rect -3442 1487 -3437 2059
rect -4019 1482 -3437 1487
rect 12681 831 12783 836
rect 12681 739 12686 831
rect 12686 739 12778 831
rect 12778 739 12783 831
rect 12681 734 12783 739
rect 19140 400 19460 720
rect -5971 -213 -5622 -208
rect -5971 -552 -5966 -213
rect -5966 -552 -5627 -213
rect -5627 -552 -5622 -213
rect -5971 -557 -5622 -552
rect 874 -306 952 -301
rect 874 -374 879 -306
rect 879 -374 947 -306
rect 947 -374 952 -306
rect 874 -379 952 -374
rect -1998 -1282 -1750 -1034
rect 3562 -306 3640 -301
rect 3562 -374 3567 -306
rect 3567 -374 3635 -306
rect 3635 -374 3640 -306
rect 3562 -379 3640 -374
rect 6250 -306 6328 -301
rect 6250 -374 6255 -306
rect 6255 -374 6323 -306
rect 6323 -374 6328 -306
rect 6250 -379 6328 -374
rect 8938 -306 9016 -301
rect 8938 -374 8943 -306
rect 8943 -374 9011 -306
rect 9011 -374 9016 -306
rect 8938 -379 9016 -374
rect 18142 -1110 18240 -1105
rect 18142 -1198 18147 -1110
rect 18147 -1198 18235 -1110
rect 18235 -1198 18240 -1110
rect 18142 -1203 18240 -1198
rect -3946 -2876 -3368 -2871
rect -3946 -3444 -3941 -2876
rect -3941 -3444 -3373 -2876
rect -3373 -3444 -3368 -2876
rect -3946 -3449 -3368 -3444
rect 3983 -2482 4393 -2477
rect 3983 -2882 3988 -2482
rect 3988 -2882 4388 -2482
rect 4388 -2882 4393 -2482
rect 3983 -2887 4393 -2882
rect 40398 -2636 40468 -2566
rect -1220 -5020 -810 -5015
rect -1220 -5420 -1215 -5020
rect -1215 -5420 -815 -5020
rect -815 -5420 -810 -5020
rect -1220 -5425 -810 -5420
rect -6018 -7150 -5622 -7145
rect -6018 -7536 -6013 -7150
rect -6013 -7536 -5627 -7150
rect -5627 -7536 -5622 -7150
rect -6018 -7541 -5622 -7536
rect -3946 -16876 -3368 -16871
rect -3946 -17444 -3941 -16876
rect -3941 -17444 -3373 -16876
rect -3373 -17444 -3368 -16876
rect -3946 -17449 -3368 -17444
rect 3983 -16482 4393 -16477
rect 3983 -16882 4080 -16482
rect 4080 -16882 4388 -16482
rect 4388 -16882 4393 -16482
rect 3983 -16887 4393 -16882
rect -1220 -19020 -810 -19015
rect -1220 -19420 -1215 -19020
rect -1215 -19420 -815 -19020
rect -815 -19420 -810 -19020
rect -1220 -19425 -810 -19420
rect -6018 -21150 -5622 -21145
rect -6018 -21536 -6013 -21150
rect -6013 -21536 -5627 -21150
rect -5627 -21536 -5622 -21150
rect -6018 -21541 -5622 -21536
rect 42446 -12036 42514 -12032
rect 42446 -12096 42450 -12036
rect 42450 -12096 42510 -12036
rect 42510 -12096 42514 -12036
rect 42446 -12100 42514 -12096
rect -3946 -30876 -3368 -30871
rect -3946 -31444 -3941 -30876
rect -3941 -31444 -3373 -30876
rect -3373 -31444 -3368 -30876
rect -3946 -31449 -3368 -31444
rect 3983 -30482 4393 -30477
rect 3983 -30882 3988 -30482
rect 3988 -30882 4388 -30482
rect 4388 -30882 4393 -30482
rect 3983 -30887 4393 -30882
rect -1220 -33020 -810 -33015
rect -1220 -33420 -1215 -33020
rect -1215 -33420 -815 -33020
rect -815 -33420 -810 -33020
rect -1220 -33425 -810 -33420
rect -6018 -35150 -5622 -35145
rect -6018 -35536 -6013 -35150
rect -6013 -35536 -5627 -35150
rect -5627 -35536 -5622 -35150
rect -6018 -35541 -5622 -35536
rect -3946 -44876 -3368 -44871
rect -3946 -45444 -3941 -44876
rect -3941 -45444 -3373 -44876
rect -3373 -45444 -3368 -44876
rect -3946 -45449 -3368 -45444
rect 3983 -44482 4393 -44477
rect 3983 -44882 3988 -44482
rect 3988 -44882 4388 -44482
rect 4388 -44882 4393 -44482
rect 3983 -44887 4393 -44882
rect -1220 -47020 -810 -47015
rect -1220 -47420 -1215 -47020
rect -1215 -47420 -815 -47020
rect -815 -47420 -810 -47020
rect -1220 -47425 -810 -47420
rect -6018 -49150 -5622 -49145
rect -6018 -49536 -6013 -49150
rect -6013 -49536 -5627 -49150
rect -5627 -49536 -5622 -49150
rect -6018 -49541 -5622 -49536
<< metal4 >>
rect -4072 2065 -3400 2092
rect -6253 -208 -5211 2025
rect -4072 1481 -4020 2065
rect -3436 1481 -3400 2065
rect -4072 1429 -3400 1481
rect 12540 945 12928 983
rect 12540 625 12572 945
rect 12892 625 12928 945
rect 12540 586 12928 625
rect 19038 720 19500 784
rect 19038 400 19140 720
rect 19460 400 19500 720
rect 19038 337 19500 400
rect -6253 -557 -5971 -208
rect -5622 -557 -5211 -208
rect 868 -301 958 -295
rect 868 -379 874 -301
rect 952 -306 958 -301
rect 3556 -301 3646 -295
rect 3556 -306 3562 -301
rect 952 -374 3562 -306
rect 952 -379 958 -374
rect 868 -385 958 -379
rect 3556 -379 3562 -374
rect 3640 -306 3646 -301
rect 6244 -301 6334 -295
rect 6244 -306 6250 -301
rect 3640 -374 6250 -306
rect 3640 -379 3646 -374
rect 3556 -385 3646 -379
rect 6244 -379 6250 -374
rect 6328 -306 6334 -301
rect 8932 -301 9022 -295
rect 8932 -306 8938 -301
rect 6328 -374 8938 -306
rect 6328 -379 6334 -374
rect 6244 -385 6334 -379
rect 8932 -379 8938 -374
rect 9016 -306 9022 -301
rect 9016 -374 12252 -306
rect 9016 -379 9022 -374
rect 8932 -385 9022 -379
rect -6253 -7145 -5211 -557
rect -2070 -998 -1654 -946
rect -2070 -1318 -2034 -998
rect -1714 -1318 -1654 -998
rect -2070 -1372 -1654 -1318
rect 12184 -2074 12252 -374
rect 17925 -994 18390 -929
rect 17925 -1314 18031 -994
rect 18351 -1314 18390 -994
rect 17925 -1367 18390 -1314
rect 12184 -2142 17212 -2074
rect 3976 -2477 4399 -2470
rect -4155 -2870 -3272 -2759
rect -4155 -3450 -3947 -2870
rect -3367 -3450 -3272 -2870
rect 3976 -2887 3983 -2477
rect 4393 -2887 4399 -2477
rect 40397 -2566 40469 -2565
rect 40397 -2636 40398 -2566
rect 40468 -2636 42515 -2566
rect 40397 -2637 40469 -2636
rect 3976 -3204 4399 -2887
rect -4155 -3608 -3272 -3450
rect -1245 -5014 -785 -4990
rect -1245 -5426 -1221 -5014
rect -809 -5426 -785 -5014
rect -1245 -5450 -785 -5426
rect -6253 -7541 -6018 -7145
rect -5622 -7541 -5211 -7145
rect -6253 -21145 -5211 -7541
rect 42445 -12016 42515 -2636
rect 42425 -12032 42537 -12016
rect 42425 -12100 42446 -12032
rect 42514 -12100 42537 -12032
rect 42425 -12114 42537 -12100
rect 3976 -16477 4399 -16470
rect -4155 -16870 -3272 -16759
rect -4155 -17450 -3947 -16870
rect -3367 -17450 -3272 -16870
rect 3976 -16887 3983 -16477
rect 4393 -16887 4399 -16477
rect 3976 -17204 4399 -16887
rect -4155 -17608 -3272 -17450
rect -1245 -19014 -785 -18990
rect -1245 -19426 -1221 -19014
rect -809 -19426 -785 -19014
rect -1245 -19450 -785 -19426
rect -6253 -21541 -6018 -21145
rect -5622 -21541 -5211 -21145
rect -6253 -35145 -5211 -21541
rect 3976 -30477 4399 -30470
rect -4155 -30870 -3272 -30759
rect -4155 -31450 -3947 -30870
rect -3367 -31450 -3272 -30870
rect 3976 -30887 3983 -30477
rect 4393 -30887 4399 -30477
rect 3976 -31204 4399 -30887
rect -4155 -31608 -3272 -31450
rect -1245 -33014 -785 -32990
rect -1245 -33426 -1221 -33014
rect -809 -33426 -785 -33014
rect -1245 -33450 -785 -33426
rect -6253 -35541 -6018 -35145
rect -5622 -35541 -5211 -35145
rect -6253 -49145 -5211 -35541
rect 3976 -44477 4399 -44470
rect -4155 -44870 -3272 -44759
rect -4155 -45450 -3947 -44870
rect -3367 -45450 -3272 -44870
rect 3976 -44887 3983 -44477
rect 4393 -44887 4399 -44477
rect 3976 -45204 4399 -44887
rect -4155 -45608 -3272 -45450
rect -1245 -47014 -785 -46990
rect -1245 -47426 -1221 -47014
rect -809 -47426 -785 -47014
rect -1245 -47450 -785 -47426
rect -6253 -49541 -6018 -49145
rect -5622 -49541 -5211 -49145
rect -6253 -57972 -5211 -49541
<< via4 >>
rect -4020 2064 -3436 2065
rect -4020 1482 -4019 2064
rect -4019 1482 -3437 2064
rect -3437 1482 -3436 2064
rect -4020 1481 -3436 1482
rect 12572 836 12892 945
rect 12572 734 12681 836
rect 12681 734 12783 836
rect 12783 734 12892 836
rect 12572 625 12892 734
rect 19140 400 19460 720
rect -2034 -1034 -1714 -998
rect -2034 -1282 -1998 -1034
rect -1998 -1282 -1750 -1034
rect -1750 -1282 -1714 -1034
rect -2034 -1318 -1714 -1282
rect 18031 -1105 18351 -994
rect 18031 -1203 18142 -1105
rect 18142 -1203 18240 -1105
rect 18240 -1203 18351 -1105
rect 18031 -1314 18351 -1203
rect -3947 -2871 -3367 -2870
rect -3947 -3449 -3946 -2871
rect -3946 -3449 -3368 -2871
rect -3368 -3449 -3367 -2871
rect -3947 -3450 -3367 -3449
rect -1221 -5015 -809 -5014
rect -1221 -5425 -1220 -5015
rect -1220 -5425 -810 -5015
rect -810 -5425 -809 -5015
rect -1221 -5426 -809 -5425
rect -3947 -16871 -3367 -16870
rect -3947 -17449 -3946 -16871
rect -3946 -17449 -3368 -16871
rect -3368 -17449 -3367 -16871
rect -3947 -17450 -3367 -17449
rect -1221 -19015 -809 -19014
rect -1221 -19425 -1220 -19015
rect -1220 -19425 -810 -19015
rect -810 -19425 -809 -19015
rect -1221 -19426 -809 -19425
rect -3947 -30871 -3367 -30870
rect -3947 -31449 -3946 -30871
rect -3946 -31449 -3368 -30871
rect -3368 -31449 -3367 -30871
rect -3947 -31450 -3367 -31449
rect -1221 -33015 -809 -33014
rect -1221 -33425 -1220 -33015
rect -1220 -33425 -810 -33015
rect -810 -33425 -809 -33015
rect -1221 -33426 -809 -33425
rect -3947 -44871 -3367 -44870
rect -3947 -45449 -3946 -44871
rect -3946 -45449 -3368 -44871
rect -3368 -45449 -3367 -44871
rect -3947 -45450 -3367 -45449
rect -1221 -47015 -809 -47014
rect -1221 -47425 -1220 -47015
rect -1220 -47425 -810 -47015
rect -810 -47425 -809 -47015
rect -1221 -47426 -809 -47425
<< metal5 >>
rect -4233 2065 -3191 2189
rect -4233 1481 -4020 2065
rect -3436 1481 -3191 2065
rect -4233 -2870 -3191 1481
rect 12459 945 13029 1132
rect 12459 625 12572 945
rect 12892 625 13029 945
rect 12459 557 13029 625
rect 19038 720 19500 784
rect 19038 400 19140 720
rect 19460 400 19500 720
rect 19038 337 19500 400
rect -2070 -998 -1654 -946
rect -2070 -1318 -2034 -998
rect -1714 -1318 -1654 -998
rect -2070 -1372 -1654 -1318
rect 17925 -994 18390 -929
rect 17925 -1314 18031 -994
rect 18351 -1314 18390 -994
rect 17925 -1367 18390 -1314
rect -4233 -3450 -3947 -2870
rect -3367 -3450 -3191 -2870
rect -4233 -16870 -3191 -3450
rect -1245 -5014 -245 -4990
rect -1245 -5426 -1221 -5014
rect -809 -5426 -245 -5014
rect -1245 -5450 -245 -5426
rect -4233 -17450 -3947 -16870
rect -3367 -17450 -3191 -16870
rect -4233 -30870 -3191 -17450
rect -1245 -19014 -245 -18990
rect -1245 -19426 -1221 -19014
rect -809 -19426 -245 -19014
rect -1245 -19450 -245 -19426
rect -4233 -31450 -3947 -30870
rect -3367 -31450 -3191 -30870
rect -4233 -44870 -3191 -31450
rect -1245 -33014 -245 -32990
rect -1245 -33426 -1221 -33014
rect -809 -33426 -245 -33014
rect -1245 -33450 -245 -33426
rect -4233 -45450 -3947 -44870
rect -3367 -45450 -3191 -44870
rect -4233 -57808 -3191 -45450
rect -1245 -47014 -245 -46990
rect -1245 -47426 -1221 -47014
rect -809 -47426 -245 -47014
rect -1245 -47450 -245 -47426
use opamp_small  opamp_small_0
timestamp 1665942972
transform 1 0 13531 0 1 -1172
box -461 -954 4014 2020
use sky130_fd_pr__cap_mim_m3_1_L4DLLG  sky130_fd_pr__cap_mim_m3_1_L4DLLG_0
timestamp 1666553439
transform 1 0 18401 0 1 -9386
box -18947 -6300 20347 6300
use sky130_fd_pr__cap_mim_m3_1_L4DLLG  sky130_fd_pr__cap_mim_m3_1_L4DLLG_1
timestamp 1666553439
transform 1 0 18401 0 1 -23386
box -18947 -6300 20347 6300
use sky130_fd_pr__cap_mim_m3_1_L4DLLG  sky130_fd_pr__cap_mim_m3_1_L4DLLG_2
timestamp 1666553439
transform 1 0 18401 0 1 -37386
box -18947 -6300 20347 6300
use sky130_fd_pr__cap_mim_m3_1_L4DLLG  sky130_fd_pr__cap_mim_m3_1_L4DLLG_3
timestamp 1666553439
transform 1 0 18401 0 1 -51386
box -18947 -6300 20347 6300
use sky130_fd_pr__cap_mim_m3_2_L4DLLG  sky130_fd_pr__cap_mim_m3_2_L4DLLG_0
timestamp 1666553597
transform 1 0 19608 0 1 -9386
box -20156 -6300 19556 6300
use sky130_fd_pr__cap_mim_m3_2_L4DLLG  sky130_fd_pr__cap_mim_m3_2_L4DLLG_1
timestamp 1666553597
transform 1 0 19608 0 1 -23386
box -20156 -6300 19556 6300
use sky130_fd_pr__cap_mim_m3_2_L4DLLG  sky130_fd_pr__cap_mim_m3_2_L4DLLG_2
timestamp 1666553597
transform 1 0 19608 0 1 -37386
box -20156 -6300 19556 6300
use sky130_fd_pr__cap_mim_m3_2_L4DLLG  sky130_fd_pr__cap_mim_m3_2_L4DLLG_3
timestamp 1666553597
transform 1 0 19608 0 1 -51386
box -20156 -6300 19556 6300
use sky130_fd_pr__nfet_01v8_lvt_9G3FLA  sky130_fd_pr__nfet_01v8_lvt_9G3FLA_0
timestamp 1666638433
transform 1 0 2861 0 1 -6451
box -647 -310 647 310
use sky130_fd_pr__nfet_01v8_lvt_9G3FLA  sky130_fd_pr__nfet_01v8_lvt_9G3FLA_1
timestamp 1666638433
transform 1 0 2861 0 1 -20451
box -647 -310 647 310
use sky130_fd_pr__nfet_01v8_lvt_9G3FLA  sky130_fd_pr__nfet_01v8_lvt_9G3FLA_2
timestamp 1666638433
transform 1 0 2861 0 1 -34451
box -647 -310 647 310
use sky130_fd_pr__nfet_01v8_lvt_9G3FLA  sky130_fd_pr__nfet_01v8_lvt_9G3FLA_3
timestamp 1666638433
transform 1 0 2861 0 1 -48451
box -647 -310 647 310
use sky130_fd_pr__nfet_01v8_lvt_R5S7KJ  sky130_fd_pr__nfet_01v8_lvt_R5S7KJ_0
timestamp 1666638433
transform 1 0 2861 0 1 -4673
box -647 -410 647 410
use sky130_fd_pr__nfet_01v8_lvt_R5S7KJ  sky130_fd_pr__nfet_01v8_lvt_R5S7KJ_1
timestamp 1666638433
transform 1 0 2861 0 1 -18673
box -647 -410 647 410
use sky130_fd_pr__nfet_01v8_lvt_R5S7KJ  sky130_fd_pr__nfet_01v8_lvt_R5S7KJ_2
timestamp 1666638433
transform 1 0 2861 0 1 -32673
box -647 -410 647 410
use sky130_fd_pr__nfet_01v8_lvt_R5S7KJ  sky130_fd_pr__nfet_01v8_lvt_R5S7KJ_3
timestamp 1666638433
transform 1 0 2861 0 1 -46673
box -647 -410 647 410
use sky130_fd_pr__nfet_g5v0d10v5_KH736R  sky130_fd_pr__nfet_g5v0d10v5_KH736R_0
timestamp 1666639277
transform 0 1 41574 -1 0 -32259
box -6519 -658 6519 658
use sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ  sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ_0
timestamp 1666571082
transform 1 0 19258 0 1 -1557
box -278 -358 278 358
use sky130_fd_pr__pfet_01v8_lvt_C38N8W  sky130_fd_pr__pfet_01v8_lvt_C38N8W_0
timestamp 1666554250
transform 1 0 1305 0 1 -4368
box -807 -719 807 719
use sky130_fd_pr__pfet_01v8_lvt_C38N8W  sky130_fd_pr__pfet_01v8_lvt_C38N8W_1
timestamp 1666554250
transform 1 0 1305 0 1 -6060
box -807 -719 807 719
use sky130_fd_pr__pfet_01v8_lvt_C38N8W  sky130_fd_pr__pfet_01v8_lvt_C38N8W_2
timestamp 1666554250
transform 1 0 1305 0 1 -18368
box -807 -719 807 719
use sky130_fd_pr__pfet_01v8_lvt_C38N8W  sky130_fd_pr__pfet_01v8_lvt_C38N8W_3
timestamp 1666554250
transform 1 0 1305 0 1 -20060
box -807 -719 807 719
use sky130_fd_pr__pfet_01v8_lvt_C38N8W  sky130_fd_pr__pfet_01v8_lvt_C38N8W_4
timestamp 1666554250
transform 1 0 1305 0 1 -32368
box -807 -719 807 719
use sky130_fd_pr__pfet_01v8_lvt_C38N8W  sky130_fd_pr__pfet_01v8_lvt_C38N8W_5
timestamp 1666554250
transform 1 0 1305 0 1 -34060
box -807 -719 807 719
use sky130_fd_pr__pfet_01v8_lvt_C38N8W  sky130_fd_pr__pfet_01v8_lvt_C38N8W_6
timestamp 1666554250
transform 1 0 1305 0 1 -46368
box -807 -719 807 719
use sky130_fd_pr__pfet_01v8_lvt_C38N8W  sky130_fd_pr__pfet_01v8_lvt_C38N8W_7
timestamp 1666554250
transform 1 0 1305 0 1 -48060
box -807 -719 807 719
use sky130_fd_pr__pfet_g5v0d10v5_5F54F3  sky130_fd_pr__pfet_g5v0d10v5_5F54F3_0
timestamp 1666639277
transform 0 1 41591 -1 0 -18214
box -6549 -697 6549 697
use sky130_fd_pr__pfet_g5v0d10v5_AJQB7U  sky130_fd_pr__pfet_g5v0d10v5_AJQB7U_0
timestamp 1666571082
transform 1 0 19246 0 1 -708
box -308 -397 308 397
use sky130_fd_pr__res_xhigh_po_0p35_RJUBBE  sky130_fd_pr__res_xhigh_po_0p35_RJUBBE_0
timestamp 1666281362
transform 0 1 13677 -1 0 -2601
box -201 -763 201 763
use sky130_fd_pr__res_xhigh_po_0p35_RJUBBE  sky130_fd_pr__res_xhigh_po_0p35_RJUBBE_1
timestamp 1666281362
transform 0 1 12147 -1 0 -2601
box -201 -763 201 763
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1661822643
transform 1 0 678 0 1 -77
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_1
timestamp 1661822643
transform 1 0 3366 0 1 -77
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_2
timestamp 1661822643
transform 1 0 6054 0 1 -77
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_3
timestamp 1661822643
transform 1 0 8742 0 1 -77
box -38 -49 2726 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1661822643
transform 1 0 2214 0 1 -1409
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_1
timestamp 1661822643
transform 1 0 4902 0 1 -1409
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_4
timestamp 1661822643
transform 1 0 7590 0 1 -1409
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_6
timestamp 1661822643
transform 1 0 10278 0 1 -1409
box -38 -49 1670 715
use sky130_fd_sc_hs__nand3_1  sky130_fd_sc_hs__nand3_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1661822643
transform 1 0 198 0 1 -77
box -38 -49 518 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1661822643
transform 1 0 6 0 1 -77
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_1
timestamp 1661822643
transform 1 0 11584 0 1 -77
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_2
timestamp 1661822643
transform -1 0 9030 0 -1 1255
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_3
timestamp 1661822643
transform -1 0 6438 0 -1 1255
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_4
timestamp 1661822643
transform -1 0 3654 0 -1 1255
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_5
timestamp 1661822643
transform -1 0 2694 0 -1 -77
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_6
timestamp 1661822643
transform 1 0 2022 0 1 -1409
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_7
timestamp 1661822643
transform 1 0 3846 0 1 -1409
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_8
timestamp 1661822643
transform -1 0 5382 0 -1 -77
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_9
timestamp 1661822643
transform -1 0 8166 0 -1 -77
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_10
timestamp 1661822643
transform -1 0 10950 0 -1 -77
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_11
timestamp 1661822643
transform 1 0 4710 0 1 -1409
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_12
timestamp 1661822643
transform 1 0 6534 0 1 -1409
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_13
timestamp 1661822643
transform 1 0 9222 0 1 -1409
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_14
timestamp 1661822643
transform 1 0 7398 0 1 -1409
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_15
timestamp 1661822643
transform 1 0 10086 0 1 -1409
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_16
timestamp 1661822643
transform 1 0 11910 0 1 -1409
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_17
timestamp 1661822643
transform -1 0 3078 0 -1 -1409
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_18
timestamp 1661822643
transform -1 0 5766 0 -1 -1409
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_19
timestamp 1661822643
transform -1 0 8358 0 -1 -1409
box -38 -49 230 715
use sky130_fd_sc_hs__tap_2  sky130_fd_sc_hs__tap_2_20
timestamp 1661822643
transform -1 0 11046 0 -1 -1409
box -38 -49 230 715
<< labels >>
rlabel metal4 -5788 1298 -5770 1308 1 GND
port 2 n
rlabel metal2 42502 -24814 42502 -24814 1 Vout
port 3 n
rlabel metal5 18034 -954 18034 -954 1 Control
port 5 n
rlabel metal5 19228 762 19228 762 1 Power
port 6 n
rlabel metal5 -1920 -966 -1920 -966 1 Clock
port 7 n
rlabel metal5 12664 1064 12664 1066 1 Ref
port 4 n
flabel metal1 s 5574 -2075 5766 -2026 0 FreeSans 200 180 0 0 VPWR
port 1 nsew power bidirectional
<< end >>
