magic
tech sky130A
magscale 1 2
timestamp 1669945358
<< obsactive >>
rect -74 5494 6226 7172
rect -74 806 818 5494
rect 5334 806 6226 5494
rect -74 -806 6226 806
rect -74 -5494 818 -806
rect 5334 -5494 6226 -806
rect -74 -7106 6226 -5494
rect -74 -11794 818 -7106
rect 5334 -11794 6226 -7106
rect -74 -13406 6226 -11794
rect -74 -18094 818 -13406
rect 5334 -18094 6226 -13406
rect -74 -19706 6226 -18094
rect -74 -24394 818 -19706
rect 5334 -24394 6226 -19706
rect -74 -26006 6226 -24394
rect -74 -30694 818 -26006
rect 5334 -30694 6226 -26006
rect -74 -32306 6226 -30694
rect -74 -36994 818 -32306
rect 5334 -36994 6226 -32306
rect -74 -38606 6226 -36994
rect -74 -43294 818 -38606
rect 5334 -43294 6226 -38606
rect -74 -44906 6226 -43294
rect -74 -49594 818 -44906
rect 5334 -49594 6226 -44906
rect -74 -51206 6226 -49594
rect -74 -55894 818 -51206
rect 5334 -55894 6226 -51206
rect -74 -57506 6226 -55894
rect -74 -62194 818 -57506
rect 5334 -62194 6226 -57506
rect -74 -63806 6226 -62194
rect -74 -68494 818 -63806
rect 5334 -68494 6226 -63806
rect -74 -70106 6226 -68494
rect -74 -74794 818 -70106
rect 5334 -74794 6226 -70106
rect -74 -76406 6226 -74794
rect -74 -81094 818 -76406
rect 5334 -81094 6226 -76406
rect -74 -82706 6226 -81094
rect -74 -87394 818 -82706
rect 5334 -87394 6226 -82706
rect -74 -89006 6226 -87394
rect -74 -93694 818 -89006
rect 5334 -93694 6226 -89006
rect -74 -95306 6226 -93694
rect -74 -99994 818 -95306
rect 5334 -99994 6226 -95306
rect -74 -101606 6226 -99994
rect -74 -106294 818 -101606
rect 5334 -106294 6226 -101606
rect -74 -107906 6226 -106294
rect -74 -112594 818 -107906
rect 5334 -112594 6226 -107906
rect -74 -114206 6226 -112594
rect -74 -118894 818 -114206
rect 5334 -118894 6226 -114206
rect -74 -120506 6226 -118894
rect -74 -125194 818 -120506
rect 5334 -125194 6226 -120506
rect -74 -126806 6226 -125194
rect -74 -131494 818 -126806
rect 5334 -131494 6226 -126806
rect -74 -133106 6226 -131494
rect -74 -137794 818 -133106
rect 5334 -137794 6226 -133106
rect -74 -139406 6226 -137794
rect -74 -144094 818 -139406
rect 5334 -144094 6226 -139406
rect -74 -145706 6226 -144094
rect -74 -150394 818 -145706
rect 5334 -150394 6226 -145706
rect -74 -152006 6226 -150394
rect -74 -156694 818 -152006
rect 5334 -156694 6226 -152006
rect -74 -158306 6226 -156694
rect -74 -162994 818 -158306
rect 5334 -162994 6226 -158306
rect -74 -164606 6226 -162994
rect -74 -169294 818 -164606
rect 5334 -169294 6226 -164606
rect -74 -170906 6226 -169294
rect -74 -175594 818 -170906
rect 5334 -175594 6226 -170906
rect -74 -177206 6226 -175594
rect -74 -181894 818 -177206
rect 5334 -181894 6226 -177206
rect -74 -183506 6226 -181894
rect -74 -188194 818 -183506
rect 5334 -188194 6226 -183506
rect -74 -189806 6226 -188194
rect -74 -194494 818 -189806
rect 5334 -194494 6226 -189806
rect -74 -196225 6226 -194494
<< metal1 >>
rect 1176 6854 1576 6874
rect 1176 6594 1196 6854
rect 1556 6594 1576 6854
rect 1176 6274 1576 6594
rect 4575 6854 4975 6874
rect 4575 6594 4595 6854
rect 4955 6594 4975 6854
rect 4575 6274 4975 6594
rect 1176 6074 4975 6274
rect 1176 -195126 1376 6074
rect 4775 -195126 4975 6074
rect 1176 -195326 4975 -195126
rect 1176 -195646 1577 -195326
rect 1176 -195906 1197 -195646
rect 1557 -195906 1577 -195646
rect 1176 -195926 1577 -195906
rect 4576 -195646 4975 -195326
rect 4576 -195906 4596 -195646
rect 4955 -195906 4975 -195646
rect 4576 -195926 4975 -195906
<< via1 >>
rect 1196 6594 1556 6854
rect 4595 6594 4955 6854
rect 1197 -195906 1557 -195646
rect 4596 -195906 4955 -195646
<< metal2 >>
rect 2776 7133 3376 7153
rect 1176 6854 1576 6874
rect 1176 6594 1196 6854
rect 1556 6594 1576 6854
rect 1176 6574 1576 6594
rect 2776 6773 2796 7133
rect 3356 6773 3376 7133
rect 2776 6424 3376 6773
rect 4575 6854 4975 6874
rect 4575 6594 4595 6854
rect 4955 6594 4975 6854
rect 4575 6574 4975 6594
rect 894 6274 5258 6424
rect 894 -195326 1044 6274
rect 5108 -195326 5258 6274
rect 894 -195476 5258 -195326
rect 1176 -195646 1577 -195626
rect 1176 -195906 1197 -195646
rect 1557 -195906 1577 -195646
rect 1176 -195926 1577 -195906
rect 2776 -195825 3376 -195476
rect 2776 -196185 2796 -195825
rect 3356 -196185 3376 -195825
rect 4576 -195646 4975 -195626
rect 4576 -195906 4596 -195646
rect 4955 -195906 4975 -195646
rect 4576 -195926 4975 -195906
rect 2776 -196205 3376 -196185
<< via2 >>
rect 1196 6594 1556 6854
rect 2796 6773 3356 7133
rect 4595 6594 4955 6854
rect 1197 -195906 1557 -195646
rect 2796 -196185 3356 -195825
rect 4596 -195906 4955 -195646
<< metal3 >>
rect 2751 7133 3394 7173
rect 1176 6854 1576 6874
rect 1176 6594 1196 6854
rect 1556 6594 1576 6854
rect 1176 6574 1576 6594
rect 2751 6773 2796 7133
rect 3356 6773 3394 7133
rect 2751 6084 3394 6773
rect 4575 6854 4975 6874
rect 4575 6594 4595 6854
rect 4955 6594 4975 6854
rect 4575 6574 4975 6594
rect 1176 -195646 1577 -195626
rect 1176 -195906 1197 -195646
rect 1557 -195906 1577 -195646
rect 1176 -195926 1577 -195906
rect 2758 -195825 3401 -195136
rect 2758 -196185 2796 -195825
rect 3356 -196185 3401 -195825
rect 4576 -195646 4975 -195626
rect 4576 -195906 4596 -195646
rect 4955 -195906 4975 -195646
rect 4576 -195926 4975 -195906
rect 2758 -196225 3401 -196185
<< via3 >>
rect 1196 6594 1556 6854
rect 2796 6773 3356 7133
rect 4595 6594 4955 6854
rect 1197 -195906 1557 -195646
rect 2796 -196185 3356 -195825
rect 4596 -195906 4955 -195646
<< metal4 >>
rect 2776 7133 3376 7153
rect 1176 6854 1576 6874
rect 1176 6594 1196 6854
rect 1556 6594 1576 6854
rect 2776 6773 2796 7133
rect 3356 6773 3376 7133
rect 2776 6753 3376 6773
rect 4575 6854 4975 6874
rect 1176 6108 1576 6594
rect 4575 6594 4595 6854
rect 4955 6594 4975 6854
rect 4575 6108 4975 6594
rect 1176 -195646 1577 -195160
rect 1176 -195906 1197 -195646
rect 1557 -195906 1577 -195646
rect 4576 -195646 4975 -195160
rect 1176 -195926 1577 -195906
rect 2776 -195825 3376 -195805
rect 2776 -196185 2796 -195825
rect 3356 -196185 3376 -195825
rect 4576 -195906 4596 -195646
rect 4955 -195906 4975 -195646
rect 4576 -195926 4975 -195906
rect 2776 -196205 3376 -196185
<< via4 >>
rect 2796 6773 3356 7133
rect 2796 -196185 3356 -195825
<< metal5 >>
rect 2751 7133 3394 7173
rect 2751 6773 2796 7133
rect 3356 6773 3394 7133
rect 2751 6084 3394 6773
rect 2758 -195825 3401 -195136
rect 2758 -196185 2796 -195825
rect 3356 -196185 3401 -195825
rect 2758 -196225 3401 -196185
use sky130_fd_pr__cap_mim_m3_1_U59KTN  sky130_fd_pr__cap_mim_m3_1_U59KTN_0
timestamp 1667066906
transform 1 0 3126 0 1 -94526
box -3200 -100800 3100 100800
use sky130_fd_pr__cap_mim_m3_2_U59KTN  sky130_fd_pr__cap_mim_m3_2_U59KTN_0
timestamp 1667067748
transform 1 0 3327 0 1 -94526
box -3401 -100800 2899 100800
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_0
timestamp 1669944869
transform 0 1 3076 -1 0 3150
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_1
timestamp 1669944869
transform 0 1 3076 -1 0 -3150
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_2
timestamp 1669944869
transform 0 1 3076 -1 0 -9450
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_3
timestamp 1669944869
transform 0 1 3076 -1 0 -15750
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_4
timestamp 1669944869
transform 0 1 3076 -1 0 -22050
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_5
timestamp 1669944869
transform 0 1 3076 -1 0 -28350
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_6
timestamp 1669944869
transform 0 1 3076 -1 0 -34650
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_7
timestamp 1669944869
transform 0 1 3076 -1 0 -40950
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_8
timestamp 1669944869
transform 0 1 3076 -1 0 -47250
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_9
timestamp 1669944869
transform 0 1 3076 -1 0 -53550
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_10
timestamp 1669944869
transform 0 1 3076 -1 0 -59850
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_11
timestamp 1669944869
transform 0 1 3076 -1 0 -66150
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_12
timestamp 1669944869
transform 0 1 3076 -1 0 -72450
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_13
timestamp 1669944869
transform 0 1 3076 -1 0 -78750
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_14
timestamp 1669944869
transform 0 1 3076 -1 0 -85050
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_15
timestamp 1669944869
transform 0 1 3076 -1 0 -91350
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_16
timestamp 1669944869
transform 0 1 3076 -1 0 -97650
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_17
timestamp 1669944869
transform 0 1 3076 -1 0 -103950
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_18
timestamp 1669944869
transform 0 1 3076 -1 0 -110250
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_19
timestamp 1669944869
transform 0 1 3076 -1 0 -116550
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_20
timestamp 1669944869
transform 0 1 3076 -1 0 -122850
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_21
timestamp 1669944869
transform 0 1 3076 -1 0 -129150
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_22
timestamp 1669944869
transform 0 1 3076 -1 0 -135450
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_23
timestamp 1669944869
transform 0 1 3076 -1 0 -141750
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_24
timestamp 1669944869
transform 0 1 3076 -1 0 -148050
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_25
timestamp 1669944869
transform 0 1 3076 -1 0 -154350
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_26
timestamp 1669944869
transform 0 1 3076 -1 0 -160650
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_27
timestamp 1669944869
transform 0 1 3076 -1 0 -166950
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_28
timestamp 1669944869
transform 0 1 3076 -1 0 -173250
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_29
timestamp 1669944869
transform 0 1 3076 -1 0 -179550
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_30
timestamp 1669944869
transform 0 1 3076 -1 0 -185850
box -2344 -2258 2344 2258
use sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ  sky130_fd_pr__nfet_g5v0d10v5_9KQQSQ_31
timestamp 1669944869
transform 0 1 3076 -1 0 -192150
box -2344 -2258 2344 2258
<< end >>
