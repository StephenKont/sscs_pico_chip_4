magic
tech sky130A
magscale 1 2
timestamp 1666045574
<< pwell >>
rect -201 -709 201 709
<< psubdiff >>
rect -165 639 -69 673
rect 69 639 165 673
rect -165 577 -131 639
rect 131 577 165 639
rect -165 -639 -131 -577
rect 131 -639 165 -577
rect -165 -673 -69 -639
rect 69 -673 165 -639
<< psubdiffcont >>
rect -69 639 69 673
rect -165 -577 -131 577
rect 131 -577 165 577
rect -69 -673 69 -639
<< xpolycontact >>
rect -35 111 35 543
rect -35 -543 35 -111
<< xpolyres >>
rect -35 -111 35 111
<< locali >>
rect -165 639 -69 673
rect 69 639 165 673
rect -165 577 -131 639
rect 131 577 165 639
rect -165 -639 -131 -577
rect 131 -639 165 -577
rect -165 -673 -69 -639
rect 69 -673 165 -639
<< viali >>
rect -19 128 19 525
rect -19 -525 19 -128
<< metal1 >>
rect -25 525 25 537
rect -25 128 -19 525
rect 19 128 25 525
rect -25 116 25 128
rect -25 -128 25 -116
rect -25 -525 -19 -128
rect 19 -525 25 -128
rect -25 -537 25 -525
<< res0p35 >>
rect -37 -113 37 113
<< properties >>
string FIXED_BBOX -148 -656 148 656
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.11 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 7.418k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
