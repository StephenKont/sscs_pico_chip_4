magic
tech sky130A
timestamp 1667515743
<< metal1 >>
rect -54525 36953 1475 37504
rect -54525 28169 -54057 36953
rect -50403 36856 1475 36953
rect -50403 28474 -5940 36856
rect 832 28474 1475 36856
rect -50403 28169 1475 28474
rect -54525 27504 1475 28169
rect 21974 36943 86474 37506
rect 21974 36811 82389 36943
rect 21974 28165 23071 36811
rect 29008 28165 82389 36811
rect 21974 28159 82389 28165
rect 86006 28159 86474 36943
rect 21974 27506 86474 28159
<< via1 >>
rect -54057 28169 -50403 36953
rect -5940 28474 832 36856
rect 23071 28165 29008 36811
rect 82389 28159 86006 36943
<< metal2 >>
rect -54525 36953 1475 37504
rect -54525 28169 -54057 36953
rect -50403 36856 1475 36953
rect -50403 28474 -5940 36856
rect 832 28474 1475 36856
rect -50403 28169 1475 28474
rect -54525 27504 1475 28169
rect 21974 36943 86474 37506
rect 21974 36811 82389 36943
rect 21974 28165 23071 36811
rect 29008 28165 82389 36811
rect 21974 28159 82389 28165
rect 86006 28159 86474 36943
rect 21974 27506 86474 28159
<< via2 >>
rect -54057 28169 -50403 36953
rect -5940 28474 832 36856
rect 23071 28165 29008 36811
rect 82389 28159 86006 36943
<< metal3 >>
rect -49026 83505 72474 91505
rect -54525 36953 -49525 37504
rect -54525 28169 -54057 36953
rect -50403 28169 -49525 36953
rect -54525 27504 -49525 28169
rect -49026 -32495 -41026 83505
rect -40526 75005 63974 83005
rect -40526 -23995 -32526 75005
rect -32026 66505 55474 74505
rect -32026 -15495 -24026 66505
rect -23526 58005 46974 66005
rect -23526 -6995 -15526 58005
rect -15026 49505 38474 57505
rect -15026 1505 -7026 49505
rect -6583 36856 1474 37504
rect -6583 28474 -5940 36856
rect 832 28474 1474 36856
rect -6583 10005 1474 28474
rect 21974 36811 29974 37506
rect 21974 28165 23071 36811
rect 29008 28165 29974 36811
rect 21974 27506 29974 28165
rect 30474 10005 38474 49505
rect -6583 2005 38474 10005
rect 38974 1505 46974 58005
rect -15026 -6495 46974 1505
rect 47474 -6995 55474 66505
rect -23526 -14995 55474 -6995
rect 55974 -15495 63974 75005
rect -32026 -23495 63974 -15495
rect 64474 -23995 72474 83505
rect 81474 36943 86474 37506
rect 81474 28159 82389 36943
rect 86006 28159 86474 36943
rect 81474 27506 86474 28159
rect -40526 -31995 72474 -23995
rect 72974 21056 86474 21505
rect 72974 13886 82020 21056
rect 85894 13886 86474 21056
rect 72974 13505 86474 13886
rect 72974 -32495 80974 13505
rect -49026 -40495 80974 -32495
<< via3 >>
rect -54057 28169 -50403 36953
rect 23071 28165 29008 36811
rect 82389 28159 86006 36943
rect 82020 13886 85894 21056
<< metal4 >>
rect -49025 83505 80975 91505
rect -49025 37504 -41025 83505
rect -54525 36953 -41025 37504
rect -54525 28169 -54057 36953
rect -50403 28169 -41025 36953
rect -54525 27504 -41025 28169
rect -40526 75006 72474 83006
rect -40526 -32494 -32526 75006
rect -32026 66506 63974 74506
rect -32026 -23994 -24026 66506
rect -23526 58006 55474 66006
rect -23526 -15494 -15526 58006
rect -15026 49506 47032 57506
rect -15026 -6994 -7026 49506
rect -6526 41006 29974 49006
rect -6526 1506 1474 41006
rect 21974 36811 29974 41006
rect 21974 28165 23071 36811
rect 29008 28165 29974 36811
rect 21974 27506 29974 28165
rect 38974 1506 47032 49506
rect -6526 -6494 47032 1506
rect 47474 -6994 55474 58006
rect -15026 -14994 55474 -6994
rect 55974 -15494 63974 66506
rect -23526 -23494 63974 -15494
rect 64474 -23994 72474 75006
rect -32026 -31994 72474 -23994
rect 72975 -32494 80975 83505
rect 81474 36943 86474 37506
rect 81474 28159 82389 36943
rect 86006 28159 86474 36943
rect 81474 27506 86474 28159
rect 81474 21056 86474 21505
rect 81474 13886 82020 21056
rect 85894 13886 86474 21056
rect 81474 13505 86474 13886
rect -40526 -40494 80975 -32494
rect 72975 -40495 80975 -40494
<< via4 >>
rect -54057 28169 -50403 36953
rect 23071 28165 29008 36811
rect 82389 28159 86006 36943
rect 82020 13886 85894 21056
<< metal5 >>
rect -49025 83505 80975 91505
rect -49025 37504 -41025 83505
rect -54525 36953 -41025 37504
rect -54525 28169 -54057 36953
rect -50403 28169 -41025 36953
rect -54525 27504 -41025 28169
rect -40526 75006 72474 83006
rect -40526 -32494 -32526 75006
rect -32026 66506 63974 74506
rect -32026 -23994 -24026 66506
rect -23526 58006 55474 66006
rect -23526 -15494 -15526 58006
rect -15026 49506 47032 57506
rect -15026 -6994 -7026 49506
rect -6526 41006 29974 49006
rect -6526 1506 1474 41006
rect 21974 36811 29974 41006
rect 21974 28165 23071 36811
rect 29008 28165 29974 36811
rect 21974 27506 29974 28165
rect 38974 1506 47032 49506
rect -6526 -6494 47032 1506
rect 47474 -6994 55474 58006
rect -15026 -14994 55474 -6994
rect 55974 -15494 63974 66506
rect -23526 -23494 63974 -15494
rect 64474 -23994 72474 75006
rect -32026 -31994 72474 -23994
rect 72975 -32494 80975 83505
rect 81474 36943 86474 37506
rect 81474 28159 82389 36943
rect 86006 28159 86474 36943
rect 81474 27506 86474 28159
rect 81474 21056 86474 21505
rect 81474 13886 82020 21056
rect 85894 13886 86474 21056
rect 81474 13505 86474 13886
rect -40526 -40494 80975 -32494
rect 72975 -40495 80975 -40494
<< end >>
