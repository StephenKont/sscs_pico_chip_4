magic
tech sky130A
magscale 1 2
timestamp 1665944614
<< pwell >>
rect -307 -720 307 720
<< psubdiff >>
rect -271 650 -175 684
rect 175 650 271 684
rect -271 588 -237 650
rect 237 588 271 650
rect -271 -650 -237 -588
rect 237 -650 271 -588
rect -271 -684 -175 -650
rect 175 -684 271 -650
<< psubdiffcont >>
rect -175 650 175 684
rect -271 -588 -237 588
rect 237 -588 271 588
rect -175 -684 175 -650
<< xpolycontact >>
rect -141 122 141 554
rect -141 -554 141 -122
<< xpolyres >>
rect -141 -122 141 122
<< locali >>
rect -271 650 -175 684
rect 175 650 271 684
rect -271 588 -237 650
rect 237 588 271 650
rect -271 -650 -237 -588
rect 237 -650 271 -588
rect -271 -684 -175 -650
rect 175 -684 271 -650
<< viali >>
rect -125 139 125 536
rect -125 -536 125 -139
<< metal1 >>
rect -131 536 131 548
rect -131 139 -125 536
rect 125 139 131 536
rect -131 127 131 139
rect -131 -139 131 -127
rect -131 -536 -125 -139
rect 125 -536 131 -139
rect -131 -548 131 -536
<< res1p41 >>
rect -143 -124 143 124
<< properties >>
string FIXED_BBOX -254 -667 254 667
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.22 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 1.997k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
