magic
tech sky130A
magscale 1 2
timestamp 1665663699
<< error_p >>
rect -927 801 -865 807
rect -799 801 -737 807
rect -671 801 -609 807
rect -543 801 -481 807
rect -415 801 -353 807
rect -287 801 -225 807
rect -159 801 -97 807
rect -31 801 31 807
rect 97 801 159 807
rect 225 801 287 807
rect 353 801 415 807
rect 481 801 543 807
rect 609 801 671 807
rect 737 801 799 807
rect 865 801 927 807
rect -927 767 -915 801
rect -799 767 -787 801
rect -671 767 -659 801
rect -543 767 -531 801
rect -415 767 -403 801
rect -287 767 -275 801
rect -159 767 -147 801
rect -31 767 -19 801
rect 97 767 109 801
rect 225 767 237 801
rect 353 767 365 801
rect 481 767 493 801
rect 609 767 621 801
rect 737 767 749 801
rect 865 767 877 801
rect -927 761 -865 767
rect -799 761 -737 767
rect -671 761 -609 767
rect -543 761 -481 767
rect -415 761 -353 767
rect -287 761 -225 767
rect -159 761 -97 767
rect -31 761 31 767
rect 97 761 159 767
rect 225 761 287 767
rect 353 761 415 767
rect 481 761 543 767
rect 609 761 671 767
rect 737 761 799 767
rect 865 761 927 767
rect -927 -767 -865 -761
rect -799 -767 -737 -761
rect -671 -767 -609 -761
rect -543 -767 -481 -761
rect -415 -767 -353 -761
rect -287 -767 -225 -761
rect -159 -767 -97 -761
rect -31 -767 31 -761
rect 97 -767 159 -761
rect 225 -767 287 -761
rect 353 -767 415 -761
rect 481 -767 543 -761
rect 609 -767 671 -761
rect 737 -767 799 -761
rect 865 -767 927 -761
rect -927 -801 -915 -767
rect -799 -801 -787 -767
rect -671 -801 -659 -767
rect -543 -801 -531 -767
rect -415 -801 -403 -767
rect -287 -801 -275 -767
rect -159 -801 -147 -767
rect -31 -801 -19 -767
rect 97 -801 109 -767
rect 225 -801 237 -767
rect 353 -801 365 -767
rect 481 -801 493 -767
rect 609 -801 621 -767
rect 737 -801 749 -767
rect 865 -801 877 -767
rect -927 -807 -865 -801
rect -799 -807 -737 -801
rect -671 -807 -609 -801
rect -543 -807 -481 -801
rect -415 -807 -353 -801
rect -287 -807 -225 -801
rect -159 -807 -97 -801
rect -31 -807 31 -801
rect 97 -807 159 -801
rect 225 -807 287 -801
rect 353 -807 415 -801
rect 481 -807 543 -801
rect 609 -807 671 -801
rect 737 -807 799 -801
rect 865 -807 927 -801
<< nwell >>
rect -1127 -939 1127 939
<< pmoslvt >>
rect -931 -720 -861 720
rect -803 -720 -733 720
rect -675 -720 -605 720
rect -547 -720 -477 720
rect -419 -720 -349 720
rect -291 -720 -221 720
rect -163 -720 -93 720
rect -35 -720 35 720
rect 93 -720 163 720
rect 221 -720 291 720
rect 349 -720 419 720
rect 477 -720 547 720
rect 605 -720 675 720
rect 733 -720 803 720
rect 861 -720 931 720
<< pdiff >>
rect -989 708 -931 720
rect -989 -708 -977 708
rect -943 -708 -931 708
rect -989 -720 -931 -708
rect -861 708 -803 720
rect -861 -708 -849 708
rect -815 -708 -803 708
rect -861 -720 -803 -708
rect -733 708 -675 720
rect -733 -708 -721 708
rect -687 -708 -675 708
rect -733 -720 -675 -708
rect -605 708 -547 720
rect -605 -708 -593 708
rect -559 -708 -547 708
rect -605 -720 -547 -708
rect -477 708 -419 720
rect -477 -708 -465 708
rect -431 -708 -419 708
rect -477 -720 -419 -708
rect -349 708 -291 720
rect -349 -708 -337 708
rect -303 -708 -291 708
rect -349 -720 -291 -708
rect -221 708 -163 720
rect -221 -708 -209 708
rect -175 -708 -163 708
rect -221 -720 -163 -708
rect -93 708 -35 720
rect -93 -708 -81 708
rect -47 -708 -35 708
rect -93 -720 -35 -708
rect 35 708 93 720
rect 35 -708 47 708
rect 81 -708 93 708
rect 35 -720 93 -708
rect 163 708 221 720
rect 163 -708 175 708
rect 209 -708 221 708
rect 163 -720 221 -708
rect 291 708 349 720
rect 291 -708 303 708
rect 337 -708 349 708
rect 291 -720 349 -708
rect 419 708 477 720
rect 419 -708 431 708
rect 465 -708 477 708
rect 419 -720 477 -708
rect 547 708 605 720
rect 547 -708 559 708
rect 593 -708 605 708
rect 547 -720 605 -708
rect 675 708 733 720
rect 675 -708 687 708
rect 721 -708 733 708
rect 675 -720 733 -708
rect 803 708 861 720
rect 803 -708 815 708
rect 849 -708 861 708
rect 803 -720 861 -708
rect 931 708 989 720
rect 931 -708 943 708
rect 977 -708 989 708
rect 931 -720 989 -708
<< pdiffc >>
rect -977 -708 -943 708
rect -849 -708 -815 708
rect -721 -708 -687 708
rect -593 -708 -559 708
rect -465 -708 -431 708
rect -337 -708 -303 708
rect -209 -708 -175 708
rect -81 -708 -47 708
rect 47 -708 81 708
rect 175 -708 209 708
rect 303 -708 337 708
rect 431 -708 465 708
rect 559 -708 593 708
rect 687 -708 721 708
rect 815 -708 849 708
rect 943 -708 977 708
<< nsubdiff >>
rect -1091 869 -995 903
rect 995 869 1091 903
rect -1091 807 -1057 869
rect 1057 807 1091 869
rect -1091 -869 -1057 -807
rect 1057 -869 1091 -807
rect -1091 -903 -995 -869
rect 995 -903 1091 -869
<< nsubdiffcont >>
rect -995 869 995 903
rect -1091 -807 -1057 807
rect 1057 -807 1091 807
rect -995 -903 995 -869
<< poly >>
rect -931 801 -861 817
rect -931 767 -915 801
rect -877 767 -861 801
rect -931 720 -861 767
rect -803 801 -733 817
rect -803 767 -787 801
rect -749 767 -733 801
rect -803 720 -733 767
rect -675 801 -605 817
rect -675 767 -659 801
rect -621 767 -605 801
rect -675 720 -605 767
rect -547 801 -477 817
rect -547 767 -531 801
rect -493 767 -477 801
rect -547 720 -477 767
rect -419 801 -349 817
rect -419 767 -403 801
rect -365 767 -349 801
rect -419 720 -349 767
rect -291 801 -221 817
rect -291 767 -275 801
rect -237 767 -221 801
rect -291 720 -221 767
rect -163 801 -93 817
rect -163 767 -147 801
rect -109 767 -93 801
rect -163 720 -93 767
rect -35 801 35 817
rect -35 767 -19 801
rect 19 767 35 801
rect -35 720 35 767
rect 93 801 163 817
rect 93 767 109 801
rect 147 767 163 801
rect 93 720 163 767
rect 221 801 291 817
rect 221 767 237 801
rect 275 767 291 801
rect 221 720 291 767
rect 349 801 419 817
rect 349 767 365 801
rect 403 767 419 801
rect 349 720 419 767
rect 477 801 547 817
rect 477 767 493 801
rect 531 767 547 801
rect 477 720 547 767
rect 605 801 675 817
rect 605 767 621 801
rect 659 767 675 801
rect 605 720 675 767
rect 733 801 803 817
rect 733 767 749 801
rect 787 767 803 801
rect 733 720 803 767
rect 861 801 931 817
rect 861 767 877 801
rect 915 767 931 801
rect 861 720 931 767
rect -931 -767 -861 -720
rect -931 -801 -915 -767
rect -877 -801 -861 -767
rect -931 -817 -861 -801
rect -803 -767 -733 -720
rect -803 -801 -787 -767
rect -749 -801 -733 -767
rect -803 -817 -733 -801
rect -675 -767 -605 -720
rect -675 -801 -659 -767
rect -621 -801 -605 -767
rect -675 -817 -605 -801
rect -547 -767 -477 -720
rect -547 -801 -531 -767
rect -493 -801 -477 -767
rect -547 -817 -477 -801
rect -419 -767 -349 -720
rect -419 -801 -403 -767
rect -365 -801 -349 -767
rect -419 -817 -349 -801
rect -291 -767 -221 -720
rect -291 -801 -275 -767
rect -237 -801 -221 -767
rect -291 -817 -221 -801
rect -163 -767 -93 -720
rect -163 -801 -147 -767
rect -109 -801 -93 -767
rect -163 -817 -93 -801
rect -35 -767 35 -720
rect -35 -801 -19 -767
rect 19 -801 35 -767
rect -35 -817 35 -801
rect 93 -767 163 -720
rect 93 -801 109 -767
rect 147 -801 163 -767
rect 93 -817 163 -801
rect 221 -767 291 -720
rect 221 -801 237 -767
rect 275 -801 291 -767
rect 221 -817 291 -801
rect 349 -767 419 -720
rect 349 -801 365 -767
rect 403 -801 419 -767
rect 349 -817 419 -801
rect 477 -767 547 -720
rect 477 -801 493 -767
rect 531 -801 547 -767
rect 477 -817 547 -801
rect 605 -767 675 -720
rect 605 -801 621 -767
rect 659 -801 675 -767
rect 605 -817 675 -801
rect 733 -767 803 -720
rect 733 -801 749 -767
rect 787 -801 803 -767
rect 733 -817 803 -801
rect 861 -767 931 -720
rect 861 -801 877 -767
rect 915 -801 931 -767
rect 861 -817 931 -801
<< polycont >>
rect -915 767 -877 801
rect -787 767 -749 801
rect -659 767 -621 801
rect -531 767 -493 801
rect -403 767 -365 801
rect -275 767 -237 801
rect -147 767 -109 801
rect -19 767 19 801
rect 109 767 147 801
rect 237 767 275 801
rect 365 767 403 801
rect 493 767 531 801
rect 621 767 659 801
rect 749 767 787 801
rect 877 767 915 801
rect -915 -801 -877 -767
rect -787 -801 -749 -767
rect -659 -801 -621 -767
rect -531 -801 -493 -767
rect -403 -801 -365 -767
rect -275 -801 -237 -767
rect -147 -801 -109 -767
rect -19 -801 19 -767
rect 109 -801 147 -767
rect 237 -801 275 -767
rect 365 -801 403 -767
rect 493 -801 531 -767
rect 621 -801 659 -767
rect 749 -801 787 -767
rect 877 -801 915 -767
<< locali >>
rect -1091 869 -995 903
rect 995 869 1091 903
rect -1091 807 -1057 869
rect 1057 807 1091 869
rect -931 767 -915 801
rect -877 767 -861 801
rect -803 767 -787 801
rect -749 767 -733 801
rect -675 767 -659 801
rect -621 767 -605 801
rect -547 767 -531 801
rect -493 767 -477 801
rect -419 767 -403 801
rect -365 767 -349 801
rect -291 767 -275 801
rect -237 767 -221 801
rect -163 767 -147 801
rect -109 767 -93 801
rect -35 767 -19 801
rect 19 767 35 801
rect 93 767 109 801
rect 147 767 163 801
rect 221 767 237 801
rect 275 767 291 801
rect 349 767 365 801
rect 403 767 419 801
rect 477 767 493 801
rect 531 767 547 801
rect 605 767 621 801
rect 659 767 675 801
rect 733 767 749 801
rect 787 767 803 801
rect 861 767 877 801
rect 915 767 931 801
rect -977 708 -943 724
rect -977 -724 -943 -708
rect -849 708 -815 724
rect -849 -724 -815 -708
rect -721 708 -687 724
rect -721 -724 -687 -708
rect -593 708 -559 724
rect -593 -724 -559 -708
rect -465 708 -431 724
rect -465 -724 -431 -708
rect -337 708 -303 724
rect -337 -724 -303 -708
rect -209 708 -175 724
rect -209 -724 -175 -708
rect -81 708 -47 724
rect -81 -724 -47 -708
rect 47 708 81 724
rect 47 -724 81 -708
rect 175 708 209 724
rect 175 -724 209 -708
rect 303 708 337 724
rect 303 -724 337 -708
rect 431 708 465 724
rect 431 -724 465 -708
rect 559 708 593 724
rect 559 -724 593 -708
rect 687 708 721 724
rect 687 -724 721 -708
rect 815 708 849 724
rect 815 -724 849 -708
rect 943 708 977 724
rect 943 -724 977 -708
rect -931 -801 -915 -767
rect -877 -801 -861 -767
rect -803 -801 -787 -767
rect -749 -801 -733 -767
rect -675 -801 -659 -767
rect -621 -801 -605 -767
rect -547 -801 -531 -767
rect -493 -801 -477 -767
rect -419 -801 -403 -767
rect -365 -801 -349 -767
rect -291 -801 -275 -767
rect -237 -801 -221 -767
rect -163 -801 -147 -767
rect -109 -801 -93 -767
rect -35 -801 -19 -767
rect 19 -801 35 -767
rect 93 -801 109 -767
rect 147 -801 163 -767
rect 221 -801 237 -767
rect 275 -801 291 -767
rect 349 -801 365 -767
rect 403 -801 419 -767
rect 477 -801 493 -767
rect 531 -801 547 -767
rect 605 -801 621 -767
rect 659 -801 675 -767
rect 733 -801 749 -767
rect 787 -801 803 -767
rect 861 -801 877 -767
rect 915 -801 931 -767
rect -1091 -869 -1057 -807
rect 1057 -869 1091 -807
rect -1091 -903 -995 -869
rect 995 -903 1091 -869
<< viali >>
rect -915 767 -877 801
rect -787 767 -749 801
rect -659 767 -621 801
rect -531 767 -493 801
rect -403 767 -365 801
rect -275 767 -237 801
rect -147 767 -109 801
rect -19 767 19 801
rect 109 767 147 801
rect 237 767 275 801
rect 365 767 403 801
rect 493 767 531 801
rect 621 767 659 801
rect 749 767 787 801
rect 877 767 915 801
rect -977 -708 -943 708
rect -849 -708 -815 708
rect -721 -708 -687 708
rect -593 -708 -559 708
rect -465 -708 -431 708
rect -337 -708 -303 708
rect -209 -708 -175 708
rect -81 -708 -47 708
rect 47 -708 81 708
rect 175 -708 209 708
rect 303 -708 337 708
rect 431 -708 465 708
rect 559 -708 593 708
rect 687 -708 721 708
rect 815 -708 849 708
rect 943 -708 977 708
rect -915 -801 -877 -767
rect -787 -801 -749 -767
rect -659 -801 -621 -767
rect -531 -801 -493 -767
rect -403 -801 -365 -767
rect -275 -801 -237 -767
rect -147 -801 -109 -767
rect -19 -801 19 -767
rect 109 -801 147 -767
rect 237 -801 275 -767
rect 365 -801 403 -767
rect 493 -801 531 -767
rect 621 -801 659 -767
rect 749 -801 787 -767
rect 877 -801 915 -767
<< metal1 >>
rect -927 801 -865 807
rect -927 767 -915 801
rect -877 767 -865 801
rect -927 761 -865 767
rect -799 801 -737 807
rect -799 767 -787 801
rect -749 767 -737 801
rect -799 761 -737 767
rect -671 801 -609 807
rect -671 767 -659 801
rect -621 767 -609 801
rect -671 761 -609 767
rect -543 801 -481 807
rect -543 767 -531 801
rect -493 767 -481 801
rect -543 761 -481 767
rect -415 801 -353 807
rect -415 767 -403 801
rect -365 767 -353 801
rect -415 761 -353 767
rect -287 801 -225 807
rect -287 767 -275 801
rect -237 767 -225 801
rect -287 761 -225 767
rect -159 801 -97 807
rect -159 767 -147 801
rect -109 767 -97 801
rect -159 761 -97 767
rect -31 801 31 807
rect -31 767 -19 801
rect 19 767 31 801
rect -31 761 31 767
rect 97 801 159 807
rect 97 767 109 801
rect 147 767 159 801
rect 97 761 159 767
rect 225 801 287 807
rect 225 767 237 801
rect 275 767 287 801
rect 225 761 287 767
rect 353 801 415 807
rect 353 767 365 801
rect 403 767 415 801
rect 353 761 415 767
rect 481 801 543 807
rect 481 767 493 801
rect 531 767 543 801
rect 481 761 543 767
rect 609 801 671 807
rect 609 767 621 801
rect 659 767 671 801
rect 609 761 671 767
rect 737 801 799 807
rect 737 767 749 801
rect 787 767 799 801
rect 737 761 799 767
rect 865 801 927 807
rect 865 767 877 801
rect 915 767 927 801
rect 865 761 927 767
rect -983 708 -937 720
rect -983 -708 -977 708
rect -943 -708 -937 708
rect -983 -720 -937 -708
rect -855 708 -809 720
rect -855 -708 -849 708
rect -815 -708 -809 708
rect -855 -720 -809 -708
rect -727 708 -681 720
rect -727 -708 -721 708
rect -687 -708 -681 708
rect -727 -720 -681 -708
rect -599 708 -553 720
rect -599 -708 -593 708
rect -559 -708 -553 708
rect -599 -720 -553 -708
rect -471 708 -425 720
rect -471 -708 -465 708
rect -431 -708 -425 708
rect -471 -720 -425 -708
rect -343 708 -297 720
rect -343 -708 -337 708
rect -303 -708 -297 708
rect -343 -720 -297 -708
rect -215 708 -169 720
rect -215 -708 -209 708
rect -175 -708 -169 708
rect -215 -720 -169 -708
rect -87 708 -41 720
rect -87 -708 -81 708
rect -47 -708 -41 708
rect -87 -720 -41 -708
rect 41 708 87 720
rect 41 -708 47 708
rect 81 -708 87 708
rect 41 -720 87 -708
rect 169 708 215 720
rect 169 -708 175 708
rect 209 -708 215 708
rect 169 -720 215 -708
rect 297 708 343 720
rect 297 -708 303 708
rect 337 -708 343 708
rect 297 -720 343 -708
rect 425 708 471 720
rect 425 -708 431 708
rect 465 -708 471 708
rect 425 -720 471 -708
rect 553 708 599 720
rect 553 -708 559 708
rect 593 -708 599 708
rect 553 -720 599 -708
rect 681 708 727 720
rect 681 -708 687 708
rect 721 -708 727 708
rect 681 -720 727 -708
rect 809 708 855 720
rect 809 -708 815 708
rect 849 -708 855 708
rect 809 -720 855 -708
rect 937 708 983 720
rect 937 -708 943 708
rect 977 -708 983 708
rect 937 -720 983 -708
rect -927 -767 -865 -761
rect -927 -801 -915 -767
rect -877 -801 -865 -767
rect -927 -807 -865 -801
rect -799 -767 -737 -761
rect -799 -801 -787 -767
rect -749 -801 -737 -767
rect -799 -807 -737 -801
rect -671 -767 -609 -761
rect -671 -801 -659 -767
rect -621 -801 -609 -767
rect -671 -807 -609 -801
rect -543 -767 -481 -761
rect -543 -801 -531 -767
rect -493 -801 -481 -767
rect -543 -807 -481 -801
rect -415 -767 -353 -761
rect -415 -801 -403 -767
rect -365 -801 -353 -767
rect -415 -807 -353 -801
rect -287 -767 -225 -761
rect -287 -801 -275 -767
rect -237 -801 -225 -767
rect -287 -807 -225 -801
rect -159 -767 -97 -761
rect -159 -801 -147 -767
rect -109 -801 -97 -767
rect -159 -807 -97 -801
rect -31 -767 31 -761
rect -31 -801 -19 -767
rect 19 -801 31 -767
rect -31 -807 31 -801
rect 97 -767 159 -761
rect 97 -801 109 -767
rect 147 -801 159 -767
rect 97 -807 159 -801
rect 225 -767 287 -761
rect 225 -801 237 -767
rect 275 -801 287 -767
rect 225 -807 287 -801
rect 353 -767 415 -761
rect 353 -801 365 -767
rect 403 -801 415 -767
rect 353 -807 415 -801
rect 481 -767 543 -761
rect 481 -801 493 -767
rect 531 -801 543 -767
rect 481 -807 543 -801
rect 609 -767 671 -761
rect 609 -801 621 -767
rect 659 -801 671 -767
rect 609 -807 671 -801
rect 737 -767 799 -761
rect 737 -801 749 -767
rect 787 -801 799 -767
rect 737 -807 799 -801
rect 865 -767 927 -761
rect 865 -801 877 -767
rect 915 -801 927 -767
rect 865 -807 927 -801
<< properties >>
string FIXED_BBOX -1074 -886 1074 886
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 7.2 l 0.35 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
