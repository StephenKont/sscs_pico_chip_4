magic
tech sky130A
magscale 1 2
timestamp 1665942972
<< error_p >>
rect -125 360 -67 366
rect 67 360 125 366
rect -125 326 -113 360
rect 67 326 79 360
rect -125 320 -67 326
rect 67 320 125 326
rect -221 -326 -163 -320
rect -29 -326 29 -320
rect 163 -326 221 -320
rect -221 -360 -209 -326
rect -29 -360 -17 -326
rect 163 -360 175 -326
rect -221 -366 -163 -360
rect -29 -366 29 -360
rect 163 -366 221 -360
<< pwell >>
rect -407 -498 407 498
<< nmoslvt >>
rect -207 -288 -177 288
rect -111 -288 -81 288
rect -15 -288 15 288
rect 81 -288 111 288
rect 177 -288 207 288
<< ndiff >>
rect -269 276 -207 288
rect -269 -276 -257 276
rect -223 -276 -207 276
rect -269 -288 -207 -276
rect -177 276 -111 288
rect -177 -276 -161 276
rect -127 -276 -111 276
rect -177 -288 -111 -276
rect -81 276 -15 288
rect -81 -276 -65 276
rect -31 -276 -15 276
rect -81 -288 -15 -276
rect 15 276 81 288
rect 15 -276 31 276
rect 65 -276 81 276
rect 15 -288 81 -276
rect 111 276 177 288
rect 111 -276 127 276
rect 161 -276 177 276
rect 111 -288 177 -276
rect 207 276 269 288
rect 207 -276 223 276
rect 257 -276 269 276
rect 207 -288 269 -276
<< ndiffc >>
rect -257 -276 -223 276
rect -161 -276 -127 276
rect -65 -276 -31 276
rect 31 -276 65 276
rect 127 -276 161 276
rect 223 -276 257 276
<< psubdiff >>
rect -371 428 -275 462
rect 275 428 371 462
rect -371 366 -337 428
rect 337 366 371 428
rect -371 -428 -337 -366
rect 337 -428 371 -366
rect -371 -462 -275 -428
rect 275 -462 371 -428
<< psubdiffcont >>
rect -275 428 275 462
rect -371 -366 -337 366
rect 337 -366 371 366
rect -275 -462 275 -428
<< poly >>
rect -129 360 -63 376
rect -129 326 -113 360
rect -79 326 -63 360
rect -207 288 -177 314
rect -129 310 -63 326
rect 63 360 129 376
rect 63 326 79 360
rect 113 326 129 360
rect -111 288 -81 310
rect -15 288 15 314
rect 63 310 129 326
rect 81 288 111 310
rect 177 288 207 314
rect -207 -310 -177 -288
rect -225 -326 -159 -310
rect -111 -314 -81 -288
rect -15 -310 15 -288
rect -225 -360 -209 -326
rect -175 -360 -159 -326
rect -225 -376 -159 -360
rect -33 -326 33 -310
rect 81 -314 111 -288
rect 177 -310 207 -288
rect -33 -360 -17 -326
rect 17 -360 33 -326
rect -33 -376 33 -360
rect 159 -326 225 -310
rect 159 -360 175 -326
rect 209 -360 225 -326
rect 159 -376 225 -360
<< polycont >>
rect -113 326 -79 360
rect 79 326 113 360
rect -209 -360 -175 -326
rect -17 -360 17 -326
rect 175 -360 209 -326
<< locali >>
rect -371 428 -275 462
rect 275 428 371 462
rect -371 366 -337 428
rect 337 366 371 428
rect -129 326 -113 360
rect -79 326 -63 360
rect 63 326 79 360
rect 113 326 129 360
rect -257 276 -223 292
rect -257 -292 -223 -276
rect -161 276 -127 292
rect -161 -292 -127 -276
rect -65 276 -31 292
rect -65 -292 -31 -276
rect 31 276 65 292
rect 31 -292 65 -276
rect 127 276 161 292
rect 127 -292 161 -276
rect 223 276 257 292
rect 223 -292 257 -276
rect -225 -360 -209 -326
rect -175 -360 -159 -326
rect -33 -360 -17 -326
rect 17 -360 33 -326
rect 159 -360 175 -326
rect 209 -360 225 -326
rect -371 -428 -337 -366
rect 337 -428 371 -366
rect -371 -462 -275 -428
rect 275 -462 371 -428
<< viali >>
rect -113 326 -79 360
rect 79 326 113 360
rect -257 -276 -223 276
rect -161 -276 -127 276
rect -65 -276 -31 276
rect 31 -276 65 276
rect 127 -276 161 276
rect 223 -276 257 276
rect -209 -360 -175 -326
rect -17 -360 17 -326
rect 175 -360 209 -326
<< metal1 >>
rect -125 360 -67 366
rect -125 326 -113 360
rect -79 326 -67 360
rect -125 320 -67 326
rect 67 360 125 366
rect 67 326 79 360
rect 113 326 125 360
rect 67 320 125 326
rect -263 276 -217 288
rect -263 -276 -257 276
rect -223 -276 -217 276
rect -263 -288 -217 -276
rect -167 276 -121 288
rect -167 -276 -161 276
rect -127 -276 -121 276
rect -167 -288 -121 -276
rect -71 276 -25 288
rect -71 -276 -65 276
rect -31 -276 -25 276
rect -71 -288 -25 -276
rect 25 276 71 288
rect 25 -276 31 276
rect 65 -276 71 276
rect 25 -288 71 -276
rect 121 276 167 288
rect 121 -276 127 276
rect 161 -276 167 276
rect 121 -288 167 -276
rect 217 276 263 288
rect 217 -276 223 276
rect 257 -276 263 276
rect 217 -288 263 -276
rect -221 -326 -163 -320
rect -221 -360 -209 -326
rect -175 -360 -163 -326
rect -221 -366 -163 -360
rect -29 -326 29 -320
rect -29 -360 -17 -326
rect 17 -360 29 -326
rect -29 -366 29 -360
rect 163 -326 221 -320
rect 163 -360 175 -326
rect 209 -360 221 -326
rect 163 -366 221 -360
<< properties >>
string FIXED_BBOX -354 -445 354 445
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.88 l 0.150 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
