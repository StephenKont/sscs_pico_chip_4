magic
tech sky130A
magscale 1 2
timestamp 1664842101
<< pwell >>
rect -1779 -1753 1779 1753
<< mvnmos >>
rect -1551 1295 -1451 1495
rect -1393 1295 -1293 1495
rect -1235 1295 -1135 1495
rect -1077 1295 -977 1495
rect -919 1295 -819 1495
rect -761 1295 -661 1495
rect -603 1295 -503 1495
rect -445 1295 -345 1495
rect -287 1295 -187 1495
rect -129 1295 -29 1495
rect 29 1295 129 1495
rect 187 1295 287 1495
rect 345 1295 445 1495
rect 503 1295 603 1495
rect 661 1295 761 1495
rect 819 1295 919 1495
rect 977 1295 1077 1495
rect 1135 1295 1235 1495
rect 1293 1295 1393 1495
rect 1451 1295 1551 1495
rect -1551 985 -1451 1185
rect -1393 985 -1293 1185
rect -1235 985 -1135 1185
rect -1077 985 -977 1185
rect -919 985 -819 1185
rect -761 985 -661 1185
rect -603 985 -503 1185
rect -445 985 -345 1185
rect -287 985 -187 1185
rect -129 985 -29 1185
rect 29 985 129 1185
rect 187 985 287 1185
rect 345 985 445 1185
rect 503 985 603 1185
rect 661 985 761 1185
rect 819 985 919 1185
rect 977 985 1077 1185
rect 1135 985 1235 1185
rect 1293 985 1393 1185
rect 1451 985 1551 1185
rect -1551 675 -1451 875
rect -1393 675 -1293 875
rect -1235 675 -1135 875
rect -1077 675 -977 875
rect -919 675 -819 875
rect -761 675 -661 875
rect -603 675 -503 875
rect -445 675 -345 875
rect -287 675 -187 875
rect -129 675 -29 875
rect 29 675 129 875
rect 187 675 287 875
rect 345 675 445 875
rect 503 675 603 875
rect 661 675 761 875
rect 819 675 919 875
rect 977 675 1077 875
rect 1135 675 1235 875
rect 1293 675 1393 875
rect 1451 675 1551 875
rect -1551 365 -1451 565
rect -1393 365 -1293 565
rect -1235 365 -1135 565
rect -1077 365 -977 565
rect -919 365 -819 565
rect -761 365 -661 565
rect -603 365 -503 565
rect -445 365 -345 565
rect -287 365 -187 565
rect -129 365 -29 565
rect 29 365 129 565
rect 187 365 287 565
rect 345 365 445 565
rect 503 365 603 565
rect 661 365 761 565
rect 819 365 919 565
rect 977 365 1077 565
rect 1135 365 1235 565
rect 1293 365 1393 565
rect 1451 365 1551 565
rect -1551 55 -1451 255
rect -1393 55 -1293 255
rect -1235 55 -1135 255
rect -1077 55 -977 255
rect -919 55 -819 255
rect -761 55 -661 255
rect -603 55 -503 255
rect -445 55 -345 255
rect -287 55 -187 255
rect -129 55 -29 255
rect 29 55 129 255
rect 187 55 287 255
rect 345 55 445 255
rect 503 55 603 255
rect 661 55 761 255
rect 819 55 919 255
rect 977 55 1077 255
rect 1135 55 1235 255
rect 1293 55 1393 255
rect 1451 55 1551 255
rect -1551 -255 -1451 -55
rect -1393 -255 -1293 -55
rect -1235 -255 -1135 -55
rect -1077 -255 -977 -55
rect -919 -255 -819 -55
rect -761 -255 -661 -55
rect -603 -255 -503 -55
rect -445 -255 -345 -55
rect -287 -255 -187 -55
rect -129 -255 -29 -55
rect 29 -255 129 -55
rect 187 -255 287 -55
rect 345 -255 445 -55
rect 503 -255 603 -55
rect 661 -255 761 -55
rect 819 -255 919 -55
rect 977 -255 1077 -55
rect 1135 -255 1235 -55
rect 1293 -255 1393 -55
rect 1451 -255 1551 -55
rect -1551 -565 -1451 -365
rect -1393 -565 -1293 -365
rect -1235 -565 -1135 -365
rect -1077 -565 -977 -365
rect -919 -565 -819 -365
rect -761 -565 -661 -365
rect -603 -565 -503 -365
rect -445 -565 -345 -365
rect -287 -565 -187 -365
rect -129 -565 -29 -365
rect 29 -565 129 -365
rect 187 -565 287 -365
rect 345 -565 445 -365
rect 503 -565 603 -365
rect 661 -565 761 -365
rect 819 -565 919 -365
rect 977 -565 1077 -365
rect 1135 -565 1235 -365
rect 1293 -565 1393 -365
rect 1451 -565 1551 -365
rect -1551 -875 -1451 -675
rect -1393 -875 -1293 -675
rect -1235 -875 -1135 -675
rect -1077 -875 -977 -675
rect -919 -875 -819 -675
rect -761 -875 -661 -675
rect -603 -875 -503 -675
rect -445 -875 -345 -675
rect -287 -875 -187 -675
rect -129 -875 -29 -675
rect 29 -875 129 -675
rect 187 -875 287 -675
rect 345 -875 445 -675
rect 503 -875 603 -675
rect 661 -875 761 -675
rect 819 -875 919 -675
rect 977 -875 1077 -675
rect 1135 -875 1235 -675
rect 1293 -875 1393 -675
rect 1451 -875 1551 -675
rect -1551 -1185 -1451 -985
rect -1393 -1185 -1293 -985
rect -1235 -1185 -1135 -985
rect -1077 -1185 -977 -985
rect -919 -1185 -819 -985
rect -761 -1185 -661 -985
rect -603 -1185 -503 -985
rect -445 -1185 -345 -985
rect -287 -1185 -187 -985
rect -129 -1185 -29 -985
rect 29 -1185 129 -985
rect 187 -1185 287 -985
rect 345 -1185 445 -985
rect 503 -1185 603 -985
rect 661 -1185 761 -985
rect 819 -1185 919 -985
rect 977 -1185 1077 -985
rect 1135 -1185 1235 -985
rect 1293 -1185 1393 -985
rect 1451 -1185 1551 -985
rect -1551 -1495 -1451 -1295
rect -1393 -1495 -1293 -1295
rect -1235 -1495 -1135 -1295
rect -1077 -1495 -977 -1295
rect -919 -1495 -819 -1295
rect -761 -1495 -661 -1295
rect -603 -1495 -503 -1295
rect -445 -1495 -345 -1295
rect -287 -1495 -187 -1295
rect -129 -1495 -29 -1295
rect 29 -1495 129 -1295
rect 187 -1495 287 -1295
rect 345 -1495 445 -1295
rect 503 -1495 603 -1295
rect 661 -1495 761 -1295
rect 819 -1495 919 -1295
rect 977 -1495 1077 -1295
rect 1135 -1495 1235 -1295
rect 1293 -1495 1393 -1295
rect 1451 -1495 1551 -1295
<< mvndiff >>
rect -1609 1483 -1551 1495
rect -1609 1307 -1597 1483
rect -1563 1307 -1551 1483
rect -1609 1295 -1551 1307
rect -1451 1483 -1393 1495
rect -1451 1307 -1439 1483
rect -1405 1307 -1393 1483
rect -1451 1295 -1393 1307
rect -1293 1483 -1235 1495
rect -1293 1307 -1281 1483
rect -1247 1307 -1235 1483
rect -1293 1295 -1235 1307
rect -1135 1483 -1077 1495
rect -1135 1307 -1123 1483
rect -1089 1307 -1077 1483
rect -1135 1295 -1077 1307
rect -977 1483 -919 1495
rect -977 1307 -965 1483
rect -931 1307 -919 1483
rect -977 1295 -919 1307
rect -819 1483 -761 1495
rect -819 1307 -807 1483
rect -773 1307 -761 1483
rect -819 1295 -761 1307
rect -661 1483 -603 1495
rect -661 1307 -649 1483
rect -615 1307 -603 1483
rect -661 1295 -603 1307
rect -503 1483 -445 1495
rect -503 1307 -491 1483
rect -457 1307 -445 1483
rect -503 1295 -445 1307
rect -345 1483 -287 1495
rect -345 1307 -333 1483
rect -299 1307 -287 1483
rect -345 1295 -287 1307
rect -187 1483 -129 1495
rect -187 1307 -175 1483
rect -141 1307 -129 1483
rect -187 1295 -129 1307
rect -29 1483 29 1495
rect -29 1307 -17 1483
rect 17 1307 29 1483
rect -29 1295 29 1307
rect 129 1483 187 1495
rect 129 1307 141 1483
rect 175 1307 187 1483
rect 129 1295 187 1307
rect 287 1483 345 1495
rect 287 1307 299 1483
rect 333 1307 345 1483
rect 287 1295 345 1307
rect 445 1483 503 1495
rect 445 1307 457 1483
rect 491 1307 503 1483
rect 445 1295 503 1307
rect 603 1483 661 1495
rect 603 1307 615 1483
rect 649 1307 661 1483
rect 603 1295 661 1307
rect 761 1483 819 1495
rect 761 1307 773 1483
rect 807 1307 819 1483
rect 761 1295 819 1307
rect 919 1483 977 1495
rect 919 1307 931 1483
rect 965 1307 977 1483
rect 919 1295 977 1307
rect 1077 1483 1135 1495
rect 1077 1307 1089 1483
rect 1123 1307 1135 1483
rect 1077 1295 1135 1307
rect 1235 1483 1293 1495
rect 1235 1307 1247 1483
rect 1281 1307 1293 1483
rect 1235 1295 1293 1307
rect 1393 1483 1451 1495
rect 1393 1307 1405 1483
rect 1439 1307 1451 1483
rect 1393 1295 1451 1307
rect 1551 1483 1609 1495
rect 1551 1307 1563 1483
rect 1597 1307 1609 1483
rect 1551 1295 1609 1307
rect -1609 1173 -1551 1185
rect -1609 997 -1597 1173
rect -1563 997 -1551 1173
rect -1609 985 -1551 997
rect -1451 1173 -1393 1185
rect -1451 997 -1439 1173
rect -1405 997 -1393 1173
rect -1451 985 -1393 997
rect -1293 1173 -1235 1185
rect -1293 997 -1281 1173
rect -1247 997 -1235 1173
rect -1293 985 -1235 997
rect -1135 1173 -1077 1185
rect -1135 997 -1123 1173
rect -1089 997 -1077 1173
rect -1135 985 -1077 997
rect -977 1173 -919 1185
rect -977 997 -965 1173
rect -931 997 -919 1173
rect -977 985 -919 997
rect -819 1173 -761 1185
rect -819 997 -807 1173
rect -773 997 -761 1173
rect -819 985 -761 997
rect -661 1173 -603 1185
rect -661 997 -649 1173
rect -615 997 -603 1173
rect -661 985 -603 997
rect -503 1173 -445 1185
rect -503 997 -491 1173
rect -457 997 -445 1173
rect -503 985 -445 997
rect -345 1173 -287 1185
rect -345 997 -333 1173
rect -299 997 -287 1173
rect -345 985 -287 997
rect -187 1173 -129 1185
rect -187 997 -175 1173
rect -141 997 -129 1173
rect -187 985 -129 997
rect -29 1173 29 1185
rect -29 997 -17 1173
rect 17 997 29 1173
rect -29 985 29 997
rect 129 1173 187 1185
rect 129 997 141 1173
rect 175 997 187 1173
rect 129 985 187 997
rect 287 1173 345 1185
rect 287 997 299 1173
rect 333 997 345 1173
rect 287 985 345 997
rect 445 1173 503 1185
rect 445 997 457 1173
rect 491 997 503 1173
rect 445 985 503 997
rect 603 1173 661 1185
rect 603 997 615 1173
rect 649 997 661 1173
rect 603 985 661 997
rect 761 1173 819 1185
rect 761 997 773 1173
rect 807 997 819 1173
rect 761 985 819 997
rect 919 1173 977 1185
rect 919 997 931 1173
rect 965 997 977 1173
rect 919 985 977 997
rect 1077 1173 1135 1185
rect 1077 997 1089 1173
rect 1123 997 1135 1173
rect 1077 985 1135 997
rect 1235 1173 1293 1185
rect 1235 997 1247 1173
rect 1281 997 1293 1173
rect 1235 985 1293 997
rect 1393 1173 1451 1185
rect 1393 997 1405 1173
rect 1439 997 1451 1173
rect 1393 985 1451 997
rect 1551 1173 1609 1185
rect 1551 997 1563 1173
rect 1597 997 1609 1173
rect 1551 985 1609 997
rect -1609 863 -1551 875
rect -1609 687 -1597 863
rect -1563 687 -1551 863
rect -1609 675 -1551 687
rect -1451 863 -1393 875
rect -1451 687 -1439 863
rect -1405 687 -1393 863
rect -1451 675 -1393 687
rect -1293 863 -1235 875
rect -1293 687 -1281 863
rect -1247 687 -1235 863
rect -1293 675 -1235 687
rect -1135 863 -1077 875
rect -1135 687 -1123 863
rect -1089 687 -1077 863
rect -1135 675 -1077 687
rect -977 863 -919 875
rect -977 687 -965 863
rect -931 687 -919 863
rect -977 675 -919 687
rect -819 863 -761 875
rect -819 687 -807 863
rect -773 687 -761 863
rect -819 675 -761 687
rect -661 863 -603 875
rect -661 687 -649 863
rect -615 687 -603 863
rect -661 675 -603 687
rect -503 863 -445 875
rect -503 687 -491 863
rect -457 687 -445 863
rect -503 675 -445 687
rect -345 863 -287 875
rect -345 687 -333 863
rect -299 687 -287 863
rect -345 675 -287 687
rect -187 863 -129 875
rect -187 687 -175 863
rect -141 687 -129 863
rect -187 675 -129 687
rect -29 863 29 875
rect -29 687 -17 863
rect 17 687 29 863
rect -29 675 29 687
rect 129 863 187 875
rect 129 687 141 863
rect 175 687 187 863
rect 129 675 187 687
rect 287 863 345 875
rect 287 687 299 863
rect 333 687 345 863
rect 287 675 345 687
rect 445 863 503 875
rect 445 687 457 863
rect 491 687 503 863
rect 445 675 503 687
rect 603 863 661 875
rect 603 687 615 863
rect 649 687 661 863
rect 603 675 661 687
rect 761 863 819 875
rect 761 687 773 863
rect 807 687 819 863
rect 761 675 819 687
rect 919 863 977 875
rect 919 687 931 863
rect 965 687 977 863
rect 919 675 977 687
rect 1077 863 1135 875
rect 1077 687 1089 863
rect 1123 687 1135 863
rect 1077 675 1135 687
rect 1235 863 1293 875
rect 1235 687 1247 863
rect 1281 687 1293 863
rect 1235 675 1293 687
rect 1393 863 1451 875
rect 1393 687 1405 863
rect 1439 687 1451 863
rect 1393 675 1451 687
rect 1551 863 1609 875
rect 1551 687 1563 863
rect 1597 687 1609 863
rect 1551 675 1609 687
rect -1609 553 -1551 565
rect -1609 377 -1597 553
rect -1563 377 -1551 553
rect -1609 365 -1551 377
rect -1451 553 -1393 565
rect -1451 377 -1439 553
rect -1405 377 -1393 553
rect -1451 365 -1393 377
rect -1293 553 -1235 565
rect -1293 377 -1281 553
rect -1247 377 -1235 553
rect -1293 365 -1235 377
rect -1135 553 -1077 565
rect -1135 377 -1123 553
rect -1089 377 -1077 553
rect -1135 365 -1077 377
rect -977 553 -919 565
rect -977 377 -965 553
rect -931 377 -919 553
rect -977 365 -919 377
rect -819 553 -761 565
rect -819 377 -807 553
rect -773 377 -761 553
rect -819 365 -761 377
rect -661 553 -603 565
rect -661 377 -649 553
rect -615 377 -603 553
rect -661 365 -603 377
rect -503 553 -445 565
rect -503 377 -491 553
rect -457 377 -445 553
rect -503 365 -445 377
rect -345 553 -287 565
rect -345 377 -333 553
rect -299 377 -287 553
rect -345 365 -287 377
rect -187 553 -129 565
rect -187 377 -175 553
rect -141 377 -129 553
rect -187 365 -129 377
rect -29 553 29 565
rect -29 377 -17 553
rect 17 377 29 553
rect -29 365 29 377
rect 129 553 187 565
rect 129 377 141 553
rect 175 377 187 553
rect 129 365 187 377
rect 287 553 345 565
rect 287 377 299 553
rect 333 377 345 553
rect 287 365 345 377
rect 445 553 503 565
rect 445 377 457 553
rect 491 377 503 553
rect 445 365 503 377
rect 603 553 661 565
rect 603 377 615 553
rect 649 377 661 553
rect 603 365 661 377
rect 761 553 819 565
rect 761 377 773 553
rect 807 377 819 553
rect 761 365 819 377
rect 919 553 977 565
rect 919 377 931 553
rect 965 377 977 553
rect 919 365 977 377
rect 1077 553 1135 565
rect 1077 377 1089 553
rect 1123 377 1135 553
rect 1077 365 1135 377
rect 1235 553 1293 565
rect 1235 377 1247 553
rect 1281 377 1293 553
rect 1235 365 1293 377
rect 1393 553 1451 565
rect 1393 377 1405 553
rect 1439 377 1451 553
rect 1393 365 1451 377
rect 1551 553 1609 565
rect 1551 377 1563 553
rect 1597 377 1609 553
rect 1551 365 1609 377
rect -1609 243 -1551 255
rect -1609 67 -1597 243
rect -1563 67 -1551 243
rect -1609 55 -1551 67
rect -1451 243 -1393 255
rect -1451 67 -1439 243
rect -1405 67 -1393 243
rect -1451 55 -1393 67
rect -1293 243 -1235 255
rect -1293 67 -1281 243
rect -1247 67 -1235 243
rect -1293 55 -1235 67
rect -1135 243 -1077 255
rect -1135 67 -1123 243
rect -1089 67 -1077 243
rect -1135 55 -1077 67
rect -977 243 -919 255
rect -977 67 -965 243
rect -931 67 -919 243
rect -977 55 -919 67
rect -819 243 -761 255
rect -819 67 -807 243
rect -773 67 -761 243
rect -819 55 -761 67
rect -661 243 -603 255
rect -661 67 -649 243
rect -615 67 -603 243
rect -661 55 -603 67
rect -503 243 -445 255
rect -503 67 -491 243
rect -457 67 -445 243
rect -503 55 -445 67
rect -345 243 -287 255
rect -345 67 -333 243
rect -299 67 -287 243
rect -345 55 -287 67
rect -187 243 -129 255
rect -187 67 -175 243
rect -141 67 -129 243
rect -187 55 -129 67
rect -29 243 29 255
rect -29 67 -17 243
rect 17 67 29 243
rect -29 55 29 67
rect 129 243 187 255
rect 129 67 141 243
rect 175 67 187 243
rect 129 55 187 67
rect 287 243 345 255
rect 287 67 299 243
rect 333 67 345 243
rect 287 55 345 67
rect 445 243 503 255
rect 445 67 457 243
rect 491 67 503 243
rect 445 55 503 67
rect 603 243 661 255
rect 603 67 615 243
rect 649 67 661 243
rect 603 55 661 67
rect 761 243 819 255
rect 761 67 773 243
rect 807 67 819 243
rect 761 55 819 67
rect 919 243 977 255
rect 919 67 931 243
rect 965 67 977 243
rect 919 55 977 67
rect 1077 243 1135 255
rect 1077 67 1089 243
rect 1123 67 1135 243
rect 1077 55 1135 67
rect 1235 243 1293 255
rect 1235 67 1247 243
rect 1281 67 1293 243
rect 1235 55 1293 67
rect 1393 243 1451 255
rect 1393 67 1405 243
rect 1439 67 1451 243
rect 1393 55 1451 67
rect 1551 243 1609 255
rect 1551 67 1563 243
rect 1597 67 1609 243
rect 1551 55 1609 67
rect -1609 -67 -1551 -55
rect -1609 -243 -1597 -67
rect -1563 -243 -1551 -67
rect -1609 -255 -1551 -243
rect -1451 -67 -1393 -55
rect -1451 -243 -1439 -67
rect -1405 -243 -1393 -67
rect -1451 -255 -1393 -243
rect -1293 -67 -1235 -55
rect -1293 -243 -1281 -67
rect -1247 -243 -1235 -67
rect -1293 -255 -1235 -243
rect -1135 -67 -1077 -55
rect -1135 -243 -1123 -67
rect -1089 -243 -1077 -67
rect -1135 -255 -1077 -243
rect -977 -67 -919 -55
rect -977 -243 -965 -67
rect -931 -243 -919 -67
rect -977 -255 -919 -243
rect -819 -67 -761 -55
rect -819 -243 -807 -67
rect -773 -243 -761 -67
rect -819 -255 -761 -243
rect -661 -67 -603 -55
rect -661 -243 -649 -67
rect -615 -243 -603 -67
rect -661 -255 -603 -243
rect -503 -67 -445 -55
rect -503 -243 -491 -67
rect -457 -243 -445 -67
rect -503 -255 -445 -243
rect -345 -67 -287 -55
rect -345 -243 -333 -67
rect -299 -243 -287 -67
rect -345 -255 -287 -243
rect -187 -67 -129 -55
rect -187 -243 -175 -67
rect -141 -243 -129 -67
rect -187 -255 -129 -243
rect -29 -67 29 -55
rect -29 -243 -17 -67
rect 17 -243 29 -67
rect -29 -255 29 -243
rect 129 -67 187 -55
rect 129 -243 141 -67
rect 175 -243 187 -67
rect 129 -255 187 -243
rect 287 -67 345 -55
rect 287 -243 299 -67
rect 333 -243 345 -67
rect 287 -255 345 -243
rect 445 -67 503 -55
rect 445 -243 457 -67
rect 491 -243 503 -67
rect 445 -255 503 -243
rect 603 -67 661 -55
rect 603 -243 615 -67
rect 649 -243 661 -67
rect 603 -255 661 -243
rect 761 -67 819 -55
rect 761 -243 773 -67
rect 807 -243 819 -67
rect 761 -255 819 -243
rect 919 -67 977 -55
rect 919 -243 931 -67
rect 965 -243 977 -67
rect 919 -255 977 -243
rect 1077 -67 1135 -55
rect 1077 -243 1089 -67
rect 1123 -243 1135 -67
rect 1077 -255 1135 -243
rect 1235 -67 1293 -55
rect 1235 -243 1247 -67
rect 1281 -243 1293 -67
rect 1235 -255 1293 -243
rect 1393 -67 1451 -55
rect 1393 -243 1405 -67
rect 1439 -243 1451 -67
rect 1393 -255 1451 -243
rect 1551 -67 1609 -55
rect 1551 -243 1563 -67
rect 1597 -243 1609 -67
rect 1551 -255 1609 -243
rect -1609 -377 -1551 -365
rect -1609 -553 -1597 -377
rect -1563 -553 -1551 -377
rect -1609 -565 -1551 -553
rect -1451 -377 -1393 -365
rect -1451 -553 -1439 -377
rect -1405 -553 -1393 -377
rect -1451 -565 -1393 -553
rect -1293 -377 -1235 -365
rect -1293 -553 -1281 -377
rect -1247 -553 -1235 -377
rect -1293 -565 -1235 -553
rect -1135 -377 -1077 -365
rect -1135 -553 -1123 -377
rect -1089 -553 -1077 -377
rect -1135 -565 -1077 -553
rect -977 -377 -919 -365
rect -977 -553 -965 -377
rect -931 -553 -919 -377
rect -977 -565 -919 -553
rect -819 -377 -761 -365
rect -819 -553 -807 -377
rect -773 -553 -761 -377
rect -819 -565 -761 -553
rect -661 -377 -603 -365
rect -661 -553 -649 -377
rect -615 -553 -603 -377
rect -661 -565 -603 -553
rect -503 -377 -445 -365
rect -503 -553 -491 -377
rect -457 -553 -445 -377
rect -503 -565 -445 -553
rect -345 -377 -287 -365
rect -345 -553 -333 -377
rect -299 -553 -287 -377
rect -345 -565 -287 -553
rect -187 -377 -129 -365
rect -187 -553 -175 -377
rect -141 -553 -129 -377
rect -187 -565 -129 -553
rect -29 -377 29 -365
rect -29 -553 -17 -377
rect 17 -553 29 -377
rect -29 -565 29 -553
rect 129 -377 187 -365
rect 129 -553 141 -377
rect 175 -553 187 -377
rect 129 -565 187 -553
rect 287 -377 345 -365
rect 287 -553 299 -377
rect 333 -553 345 -377
rect 287 -565 345 -553
rect 445 -377 503 -365
rect 445 -553 457 -377
rect 491 -553 503 -377
rect 445 -565 503 -553
rect 603 -377 661 -365
rect 603 -553 615 -377
rect 649 -553 661 -377
rect 603 -565 661 -553
rect 761 -377 819 -365
rect 761 -553 773 -377
rect 807 -553 819 -377
rect 761 -565 819 -553
rect 919 -377 977 -365
rect 919 -553 931 -377
rect 965 -553 977 -377
rect 919 -565 977 -553
rect 1077 -377 1135 -365
rect 1077 -553 1089 -377
rect 1123 -553 1135 -377
rect 1077 -565 1135 -553
rect 1235 -377 1293 -365
rect 1235 -553 1247 -377
rect 1281 -553 1293 -377
rect 1235 -565 1293 -553
rect 1393 -377 1451 -365
rect 1393 -553 1405 -377
rect 1439 -553 1451 -377
rect 1393 -565 1451 -553
rect 1551 -377 1609 -365
rect 1551 -553 1563 -377
rect 1597 -553 1609 -377
rect 1551 -565 1609 -553
rect -1609 -687 -1551 -675
rect -1609 -863 -1597 -687
rect -1563 -863 -1551 -687
rect -1609 -875 -1551 -863
rect -1451 -687 -1393 -675
rect -1451 -863 -1439 -687
rect -1405 -863 -1393 -687
rect -1451 -875 -1393 -863
rect -1293 -687 -1235 -675
rect -1293 -863 -1281 -687
rect -1247 -863 -1235 -687
rect -1293 -875 -1235 -863
rect -1135 -687 -1077 -675
rect -1135 -863 -1123 -687
rect -1089 -863 -1077 -687
rect -1135 -875 -1077 -863
rect -977 -687 -919 -675
rect -977 -863 -965 -687
rect -931 -863 -919 -687
rect -977 -875 -919 -863
rect -819 -687 -761 -675
rect -819 -863 -807 -687
rect -773 -863 -761 -687
rect -819 -875 -761 -863
rect -661 -687 -603 -675
rect -661 -863 -649 -687
rect -615 -863 -603 -687
rect -661 -875 -603 -863
rect -503 -687 -445 -675
rect -503 -863 -491 -687
rect -457 -863 -445 -687
rect -503 -875 -445 -863
rect -345 -687 -287 -675
rect -345 -863 -333 -687
rect -299 -863 -287 -687
rect -345 -875 -287 -863
rect -187 -687 -129 -675
rect -187 -863 -175 -687
rect -141 -863 -129 -687
rect -187 -875 -129 -863
rect -29 -687 29 -675
rect -29 -863 -17 -687
rect 17 -863 29 -687
rect -29 -875 29 -863
rect 129 -687 187 -675
rect 129 -863 141 -687
rect 175 -863 187 -687
rect 129 -875 187 -863
rect 287 -687 345 -675
rect 287 -863 299 -687
rect 333 -863 345 -687
rect 287 -875 345 -863
rect 445 -687 503 -675
rect 445 -863 457 -687
rect 491 -863 503 -687
rect 445 -875 503 -863
rect 603 -687 661 -675
rect 603 -863 615 -687
rect 649 -863 661 -687
rect 603 -875 661 -863
rect 761 -687 819 -675
rect 761 -863 773 -687
rect 807 -863 819 -687
rect 761 -875 819 -863
rect 919 -687 977 -675
rect 919 -863 931 -687
rect 965 -863 977 -687
rect 919 -875 977 -863
rect 1077 -687 1135 -675
rect 1077 -863 1089 -687
rect 1123 -863 1135 -687
rect 1077 -875 1135 -863
rect 1235 -687 1293 -675
rect 1235 -863 1247 -687
rect 1281 -863 1293 -687
rect 1235 -875 1293 -863
rect 1393 -687 1451 -675
rect 1393 -863 1405 -687
rect 1439 -863 1451 -687
rect 1393 -875 1451 -863
rect 1551 -687 1609 -675
rect 1551 -863 1563 -687
rect 1597 -863 1609 -687
rect 1551 -875 1609 -863
rect -1609 -997 -1551 -985
rect -1609 -1173 -1597 -997
rect -1563 -1173 -1551 -997
rect -1609 -1185 -1551 -1173
rect -1451 -997 -1393 -985
rect -1451 -1173 -1439 -997
rect -1405 -1173 -1393 -997
rect -1451 -1185 -1393 -1173
rect -1293 -997 -1235 -985
rect -1293 -1173 -1281 -997
rect -1247 -1173 -1235 -997
rect -1293 -1185 -1235 -1173
rect -1135 -997 -1077 -985
rect -1135 -1173 -1123 -997
rect -1089 -1173 -1077 -997
rect -1135 -1185 -1077 -1173
rect -977 -997 -919 -985
rect -977 -1173 -965 -997
rect -931 -1173 -919 -997
rect -977 -1185 -919 -1173
rect -819 -997 -761 -985
rect -819 -1173 -807 -997
rect -773 -1173 -761 -997
rect -819 -1185 -761 -1173
rect -661 -997 -603 -985
rect -661 -1173 -649 -997
rect -615 -1173 -603 -997
rect -661 -1185 -603 -1173
rect -503 -997 -445 -985
rect -503 -1173 -491 -997
rect -457 -1173 -445 -997
rect -503 -1185 -445 -1173
rect -345 -997 -287 -985
rect -345 -1173 -333 -997
rect -299 -1173 -287 -997
rect -345 -1185 -287 -1173
rect -187 -997 -129 -985
rect -187 -1173 -175 -997
rect -141 -1173 -129 -997
rect -187 -1185 -129 -1173
rect -29 -997 29 -985
rect -29 -1173 -17 -997
rect 17 -1173 29 -997
rect -29 -1185 29 -1173
rect 129 -997 187 -985
rect 129 -1173 141 -997
rect 175 -1173 187 -997
rect 129 -1185 187 -1173
rect 287 -997 345 -985
rect 287 -1173 299 -997
rect 333 -1173 345 -997
rect 287 -1185 345 -1173
rect 445 -997 503 -985
rect 445 -1173 457 -997
rect 491 -1173 503 -997
rect 445 -1185 503 -1173
rect 603 -997 661 -985
rect 603 -1173 615 -997
rect 649 -1173 661 -997
rect 603 -1185 661 -1173
rect 761 -997 819 -985
rect 761 -1173 773 -997
rect 807 -1173 819 -997
rect 761 -1185 819 -1173
rect 919 -997 977 -985
rect 919 -1173 931 -997
rect 965 -1173 977 -997
rect 919 -1185 977 -1173
rect 1077 -997 1135 -985
rect 1077 -1173 1089 -997
rect 1123 -1173 1135 -997
rect 1077 -1185 1135 -1173
rect 1235 -997 1293 -985
rect 1235 -1173 1247 -997
rect 1281 -1173 1293 -997
rect 1235 -1185 1293 -1173
rect 1393 -997 1451 -985
rect 1393 -1173 1405 -997
rect 1439 -1173 1451 -997
rect 1393 -1185 1451 -1173
rect 1551 -997 1609 -985
rect 1551 -1173 1563 -997
rect 1597 -1173 1609 -997
rect 1551 -1185 1609 -1173
rect -1609 -1307 -1551 -1295
rect -1609 -1483 -1597 -1307
rect -1563 -1483 -1551 -1307
rect -1609 -1495 -1551 -1483
rect -1451 -1307 -1393 -1295
rect -1451 -1483 -1439 -1307
rect -1405 -1483 -1393 -1307
rect -1451 -1495 -1393 -1483
rect -1293 -1307 -1235 -1295
rect -1293 -1483 -1281 -1307
rect -1247 -1483 -1235 -1307
rect -1293 -1495 -1235 -1483
rect -1135 -1307 -1077 -1295
rect -1135 -1483 -1123 -1307
rect -1089 -1483 -1077 -1307
rect -1135 -1495 -1077 -1483
rect -977 -1307 -919 -1295
rect -977 -1483 -965 -1307
rect -931 -1483 -919 -1307
rect -977 -1495 -919 -1483
rect -819 -1307 -761 -1295
rect -819 -1483 -807 -1307
rect -773 -1483 -761 -1307
rect -819 -1495 -761 -1483
rect -661 -1307 -603 -1295
rect -661 -1483 -649 -1307
rect -615 -1483 -603 -1307
rect -661 -1495 -603 -1483
rect -503 -1307 -445 -1295
rect -503 -1483 -491 -1307
rect -457 -1483 -445 -1307
rect -503 -1495 -445 -1483
rect -345 -1307 -287 -1295
rect -345 -1483 -333 -1307
rect -299 -1483 -287 -1307
rect -345 -1495 -287 -1483
rect -187 -1307 -129 -1295
rect -187 -1483 -175 -1307
rect -141 -1483 -129 -1307
rect -187 -1495 -129 -1483
rect -29 -1307 29 -1295
rect -29 -1483 -17 -1307
rect 17 -1483 29 -1307
rect -29 -1495 29 -1483
rect 129 -1307 187 -1295
rect 129 -1483 141 -1307
rect 175 -1483 187 -1307
rect 129 -1495 187 -1483
rect 287 -1307 345 -1295
rect 287 -1483 299 -1307
rect 333 -1483 345 -1307
rect 287 -1495 345 -1483
rect 445 -1307 503 -1295
rect 445 -1483 457 -1307
rect 491 -1483 503 -1307
rect 445 -1495 503 -1483
rect 603 -1307 661 -1295
rect 603 -1483 615 -1307
rect 649 -1483 661 -1307
rect 603 -1495 661 -1483
rect 761 -1307 819 -1295
rect 761 -1483 773 -1307
rect 807 -1483 819 -1307
rect 761 -1495 819 -1483
rect 919 -1307 977 -1295
rect 919 -1483 931 -1307
rect 965 -1483 977 -1307
rect 919 -1495 977 -1483
rect 1077 -1307 1135 -1295
rect 1077 -1483 1089 -1307
rect 1123 -1483 1135 -1307
rect 1077 -1495 1135 -1483
rect 1235 -1307 1293 -1295
rect 1235 -1483 1247 -1307
rect 1281 -1483 1293 -1307
rect 1235 -1495 1293 -1483
rect 1393 -1307 1451 -1295
rect 1393 -1483 1405 -1307
rect 1439 -1483 1451 -1307
rect 1393 -1495 1451 -1483
rect 1551 -1307 1609 -1295
rect 1551 -1483 1563 -1307
rect 1597 -1483 1609 -1307
rect 1551 -1495 1609 -1483
<< mvndiffc >>
rect -1597 1307 -1563 1483
rect -1439 1307 -1405 1483
rect -1281 1307 -1247 1483
rect -1123 1307 -1089 1483
rect -965 1307 -931 1483
rect -807 1307 -773 1483
rect -649 1307 -615 1483
rect -491 1307 -457 1483
rect -333 1307 -299 1483
rect -175 1307 -141 1483
rect -17 1307 17 1483
rect 141 1307 175 1483
rect 299 1307 333 1483
rect 457 1307 491 1483
rect 615 1307 649 1483
rect 773 1307 807 1483
rect 931 1307 965 1483
rect 1089 1307 1123 1483
rect 1247 1307 1281 1483
rect 1405 1307 1439 1483
rect 1563 1307 1597 1483
rect -1597 997 -1563 1173
rect -1439 997 -1405 1173
rect -1281 997 -1247 1173
rect -1123 997 -1089 1173
rect -965 997 -931 1173
rect -807 997 -773 1173
rect -649 997 -615 1173
rect -491 997 -457 1173
rect -333 997 -299 1173
rect -175 997 -141 1173
rect -17 997 17 1173
rect 141 997 175 1173
rect 299 997 333 1173
rect 457 997 491 1173
rect 615 997 649 1173
rect 773 997 807 1173
rect 931 997 965 1173
rect 1089 997 1123 1173
rect 1247 997 1281 1173
rect 1405 997 1439 1173
rect 1563 997 1597 1173
rect -1597 687 -1563 863
rect -1439 687 -1405 863
rect -1281 687 -1247 863
rect -1123 687 -1089 863
rect -965 687 -931 863
rect -807 687 -773 863
rect -649 687 -615 863
rect -491 687 -457 863
rect -333 687 -299 863
rect -175 687 -141 863
rect -17 687 17 863
rect 141 687 175 863
rect 299 687 333 863
rect 457 687 491 863
rect 615 687 649 863
rect 773 687 807 863
rect 931 687 965 863
rect 1089 687 1123 863
rect 1247 687 1281 863
rect 1405 687 1439 863
rect 1563 687 1597 863
rect -1597 377 -1563 553
rect -1439 377 -1405 553
rect -1281 377 -1247 553
rect -1123 377 -1089 553
rect -965 377 -931 553
rect -807 377 -773 553
rect -649 377 -615 553
rect -491 377 -457 553
rect -333 377 -299 553
rect -175 377 -141 553
rect -17 377 17 553
rect 141 377 175 553
rect 299 377 333 553
rect 457 377 491 553
rect 615 377 649 553
rect 773 377 807 553
rect 931 377 965 553
rect 1089 377 1123 553
rect 1247 377 1281 553
rect 1405 377 1439 553
rect 1563 377 1597 553
rect -1597 67 -1563 243
rect -1439 67 -1405 243
rect -1281 67 -1247 243
rect -1123 67 -1089 243
rect -965 67 -931 243
rect -807 67 -773 243
rect -649 67 -615 243
rect -491 67 -457 243
rect -333 67 -299 243
rect -175 67 -141 243
rect -17 67 17 243
rect 141 67 175 243
rect 299 67 333 243
rect 457 67 491 243
rect 615 67 649 243
rect 773 67 807 243
rect 931 67 965 243
rect 1089 67 1123 243
rect 1247 67 1281 243
rect 1405 67 1439 243
rect 1563 67 1597 243
rect -1597 -243 -1563 -67
rect -1439 -243 -1405 -67
rect -1281 -243 -1247 -67
rect -1123 -243 -1089 -67
rect -965 -243 -931 -67
rect -807 -243 -773 -67
rect -649 -243 -615 -67
rect -491 -243 -457 -67
rect -333 -243 -299 -67
rect -175 -243 -141 -67
rect -17 -243 17 -67
rect 141 -243 175 -67
rect 299 -243 333 -67
rect 457 -243 491 -67
rect 615 -243 649 -67
rect 773 -243 807 -67
rect 931 -243 965 -67
rect 1089 -243 1123 -67
rect 1247 -243 1281 -67
rect 1405 -243 1439 -67
rect 1563 -243 1597 -67
rect -1597 -553 -1563 -377
rect -1439 -553 -1405 -377
rect -1281 -553 -1247 -377
rect -1123 -553 -1089 -377
rect -965 -553 -931 -377
rect -807 -553 -773 -377
rect -649 -553 -615 -377
rect -491 -553 -457 -377
rect -333 -553 -299 -377
rect -175 -553 -141 -377
rect -17 -553 17 -377
rect 141 -553 175 -377
rect 299 -553 333 -377
rect 457 -553 491 -377
rect 615 -553 649 -377
rect 773 -553 807 -377
rect 931 -553 965 -377
rect 1089 -553 1123 -377
rect 1247 -553 1281 -377
rect 1405 -553 1439 -377
rect 1563 -553 1597 -377
rect -1597 -863 -1563 -687
rect -1439 -863 -1405 -687
rect -1281 -863 -1247 -687
rect -1123 -863 -1089 -687
rect -965 -863 -931 -687
rect -807 -863 -773 -687
rect -649 -863 -615 -687
rect -491 -863 -457 -687
rect -333 -863 -299 -687
rect -175 -863 -141 -687
rect -17 -863 17 -687
rect 141 -863 175 -687
rect 299 -863 333 -687
rect 457 -863 491 -687
rect 615 -863 649 -687
rect 773 -863 807 -687
rect 931 -863 965 -687
rect 1089 -863 1123 -687
rect 1247 -863 1281 -687
rect 1405 -863 1439 -687
rect 1563 -863 1597 -687
rect -1597 -1173 -1563 -997
rect -1439 -1173 -1405 -997
rect -1281 -1173 -1247 -997
rect -1123 -1173 -1089 -997
rect -965 -1173 -931 -997
rect -807 -1173 -773 -997
rect -649 -1173 -615 -997
rect -491 -1173 -457 -997
rect -333 -1173 -299 -997
rect -175 -1173 -141 -997
rect -17 -1173 17 -997
rect 141 -1173 175 -997
rect 299 -1173 333 -997
rect 457 -1173 491 -997
rect 615 -1173 649 -997
rect 773 -1173 807 -997
rect 931 -1173 965 -997
rect 1089 -1173 1123 -997
rect 1247 -1173 1281 -997
rect 1405 -1173 1439 -997
rect 1563 -1173 1597 -997
rect -1597 -1483 -1563 -1307
rect -1439 -1483 -1405 -1307
rect -1281 -1483 -1247 -1307
rect -1123 -1483 -1089 -1307
rect -965 -1483 -931 -1307
rect -807 -1483 -773 -1307
rect -649 -1483 -615 -1307
rect -491 -1483 -457 -1307
rect -333 -1483 -299 -1307
rect -175 -1483 -141 -1307
rect -17 -1483 17 -1307
rect 141 -1483 175 -1307
rect 299 -1483 333 -1307
rect 457 -1483 491 -1307
rect 615 -1483 649 -1307
rect 773 -1483 807 -1307
rect 931 -1483 965 -1307
rect 1089 -1483 1123 -1307
rect 1247 -1483 1281 -1307
rect 1405 -1483 1439 -1307
rect 1563 -1483 1597 -1307
<< mvpsubdiff >>
rect -1743 1705 1743 1717
rect -1743 1671 -1635 1705
rect 1635 1671 1743 1705
rect -1743 1659 1743 1671
rect -1743 1609 -1685 1659
rect -1743 -1609 -1731 1609
rect -1697 -1609 -1685 1609
rect 1685 1609 1743 1659
rect -1743 -1659 -1685 -1609
rect 1685 -1609 1697 1609
rect 1731 -1609 1743 1609
rect 1685 -1659 1743 -1609
rect -1743 -1671 1743 -1659
rect -1743 -1705 -1635 -1671
rect 1635 -1705 1743 -1671
rect -1743 -1717 1743 -1705
<< mvpsubdiffcont >>
rect -1635 1671 1635 1705
rect -1731 -1609 -1697 1609
rect 1697 -1609 1731 1609
rect -1635 -1705 1635 -1671
<< poly >>
rect -1551 1567 -1451 1583
rect -1551 1533 -1535 1567
rect -1467 1533 -1451 1567
rect -1551 1495 -1451 1533
rect -1393 1567 -1293 1583
rect -1393 1533 -1377 1567
rect -1309 1533 -1293 1567
rect -1393 1495 -1293 1533
rect -1235 1567 -1135 1583
rect -1235 1533 -1219 1567
rect -1151 1533 -1135 1567
rect -1235 1495 -1135 1533
rect -1077 1567 -977 1583
rect -1077 1533 -1061 1567
rect -993 1533 -977 1567
rect -1077 1495 -977 1533
rect -919 1567 -819 1583
rect -919 1533 -903 1567
rect -835 1533 -819 1567
rect -919 1495 -819 1533
rect -761 1567 -661 1583
rect -761 1533 -745 1567
rect -677 1533 -661 1567
rect -761 1495 -661 1533
rect -603 1567 -503 1583
rect -603 1533 -587 1567
rect -519 1533 -503 1567
rect -603 1495 -503 1533
rect -445 1567 -345 1583
rect -445 1533 -429 1567
rect -361 1533 -345 1567
rect -445 1495 -345 1533
rect -287 1567 -187 1583
rect -287 1533 -271 1567
rect -203 1533 -187 1567
rect -287 1495 -187 1533
rect -129 1567 -29 1583
rect -129 1533 -113 1567
rect -45 1533 -29 1567
rect -129 1495 -29 1533
rect 29 1567 129 1583
rect 29 1533 45 1567
rect 113 1533 129 1567
rect 29 1495 129 1533
rect 187 1567 287 1583
rect 187 1533 203 1567
rect 271 1533 287 1567
rect 187 1495 287 1533
rect 345 1567 445 1583
rect 345 1533 361 1567
rect 429 1533 445 1567
rect 345 1495 445 1533
rect 503 1567 603 1583
rect 503 1533 519 1567
rect 587 1533 603 1567
rect 503 1495 603 1533
rect 661 1567 761 1583
rect 661 1533 677 1567
rect 745 1533 761 1567
rect 661 1495 761 1533
rect 819 1567 919 1583
rect 819 1533 835 1567
rect 903 1533 919 1567
rect 819 1495 919 1533
rect 977 1567 1077 1583
rect 977 1533 993 1567
rect 1061 1533 1077 1567
rect 977 1495 1077 1533
rect 1135 1567 1235 1583
rect 1135 1533 1151 1567
rect 1219 1533 1235 1567
rect 1135 1495 1235 1533
rect 1293 1567 1393 1583
rect 1293 1533 1309 1567
rect 1377 1533 1393 1567
rect 1293 1495 1393 1533
rect 1451 1567 1551 1583
rect 1451 1533 1467 1567
rect 1535 1533 1551 1567
rect 1451 1495 1551 1533
rect -1551 1257 -1451 1295
rect -1551 1223 -1535 1257
rect -1467 1223 -1451 1257
rect -1551 1185 -1451 1223
rect -1393 1257 -1293 1295
rect -1393 1223 -1377 1257
rect -1309 1223 -1293 1257
rect -1393 1185 -1293 1223
rect -1235 1257 -1135 1295
rect -1235 1223 -1219 1257
rect -1151 1223 -1135 1257
rect -1235 1185 -1135 1223
rect -1077 1257 -977 1295
rect -1077 1223 -1061 1257
rect -993 1223 -977 1257
rect -1077 1185 -977 1223
rect -919 1257 -819 1295
rect -919 1223 -903 1257
rect -835 1223 -819 1257
rect -919 1185 -819 1223
rect -761 1257 -661 1295
rect -761 1223 -745 1257
rect -677 1223 -661 1257
rect -761 1185 -661 1223
rect -603 1257 -503 1295
rect -603 1223 -587 1257
rect -519 1223 -503 1257
rect -603 1185 -503 1223
rect -445 1257 -345 1295
rect -445 1223 -429 1257
rect -361 1223 -345 1257
rect -445 1185 -345 1223
rect -287 1257 -187 1295
rect -287 1223 -271 1257
rect -203 1223 -187 1257
rect -287 1185 -187 1223
rect -129 1257 -29 1295
rect -129 1223 -113 1257
rect -45 1223 -29 1257
rect -129 1185 -29 1223
rect 29 1257 129 1295
rect 29 1223 45 1257
rect 113 1223 129 1257
rect 29 1185 129 1223
rect 187 1257 287 1295
rect 187 1223 203 1257
rect 271 1223 287 1257
rect 187 1185 287 1223
rect 345 1257 445 1295
rect 345 1223 361 1257
rect 429 1223 445 1257
rect 345 1185 445 1223
rect 503 1257 603 1295
rect 503 1223 519 1257
rect 587 1223 603 1257
rect 503 1185 603 1223
rect 661 1257 761 1295
rect 661 1223 677 1257
rect 745 1223 761 1257
rect 661 1185 761 1223
rect 819 1257 919 1295
rect 819 1223 835 1257
rect 903 1223 919 1257
rect 819 1185 919 1223
rect 977 1257 1077 1295
rect 977 1223 993 1257
rect 1061 1223 1077 1257
rect 977 1185 1077 1223
rect 1135 1257 1235 1295
rect 1135 1223 1151 1257
rect 1219 1223 1235 1257
rect 1135 1185 1235 1223
rect 1293 1257 1393 1295
rect 1293 1223 1309 1257
rect 1377 1223 1393 1257
rect 1293 1185 1393 1223
rect 1451 1257 1551 1295
rect 1451 1223 1467 1257
rect 1535 1223 1551 1257
rect 1451 1185 1551 1223
rect -1551 947 -1451 985
rect -1551 913 -1535 947
rect -1467 913 -1451 947
rect -1551 875 -1451 913
rect -1393 947 -1293 985
rect -1393 913 -1377 947
rect -1309 913 -1293 947
rect -1393 875 -1293 913
rect -1235 947 -1135 985
rect -1235 913 -1219 947
rect -1151 913 -1135 947
rect -1235 875 -1135 913
rect -1077 947 -977 985
rect -1077 913 -1061 947
rect -993 913 -977 947
rect -1077 875 -977 913
rect -919 947 -819 985
rect -919 913 -903 947
rect -835 913 -819 947
rect -919 875 -819 913
rect -761 947 -661 985
rect -761 913 -745 947
rect -677 913 -661 947
rect -761 875 -661 913
rect -603 947 -503 985
rect -603 913 -587 947
rect -519 913 -503 947
rect -603 875 -503 913
rect -445 947 -345 985
rect -445 913 -429 947
rect -361 913 -345 947
rect -445 875 -345 913
rect -287 947 -187 985
rect -287 913 -271 947
rect -203 913 -187 947
rect -287 875 -187 913
rect -129 947 -29 985
rect -129 913 -113 947
rect -45 913 -29 947
rect -129 875 -29 913
rect 29 947 129 985
rect 29 913 45 947
rect 113 913 129 947
rect 29 875 129 913
rect 187 947 287 985
rect 187 913 203 947
rect 271 913 287 947
rect 187 875 287 913
rect 345 947 445 985
rect 345 913 361 947
rect 429 913 445 947
rect 345 875 445 913
rect 503 947 603 985
rect 503 913 519 947
rect 587 913 603 947
rect 503 875 603 913
rect 661 947 761 985
rect 661 913 677 947
rect 745 913 761 947
rect 661 875 761 913
rect 819 947 919 985
rect 819 913 835 947
rect 903 913 919 947
rect 819 875 919 913
rect 977 947 1077 985
rect 977 913 993 947
rect 1061 913 1077 947
rect 977 875 1077 913
rect 1135 947 1235 985
rect 1135 913 1151 947
rect 1219 913 1235 947
rect 1135 875 1235 913
rect 1293 947 1393 985
rect 1293 913 1309 947
rect 1377 913 1393 947
rect 1293 875 1393 913
rect 1451 947 1551 985
rect 1451 913 1467 947
rect 1535 913 1551 947
rect 1451 875 1551 913
rect -1551 637 -1451 675
rect -1551 603 -1535 637
rect -1467 603 -1451 637
rect -1551 565 -1451 603
rect -1393 637 -1293 675
rect -1393 603 -1377 637
rect -1309 603 -1293 637
rect -1393 565 -1293 603
rect -1235 637 -1135 675
rect -1235 603 -1219 637
rect -1151 603 -1135 637
rect -1235 565 -1135 603
rect -1077 637 -977 675
rect -1077 603 -1061 637
rect -993 603 -977 637
rect -1077 565 -977 603
rect -919 637 -819 675
rect -919 603 -903 637
rect -835 603 -819 637
rect -919 565 -819 603
rect -761 637 -661 675
rect -761 603 -745 637
rect -677 603 -661 637
rect -761 565 -661 603
rect -603 637 -503 675
rect -603 603 -587 637
rect -519 603 -503 637
rect -603 565 -503 603
rect -445 637 -345 675
rect -445 603 -429 637
rect -361 603 -345 637
rect -445 565 -345 603
rect -287 637 -187 675
rect -287 603 -271 637
rect -203 603 -187 637
rect -287 565 -187 603
rect -129 637 -29 675
rect -129 603 -113 637
rect -45 603 -29 637
rect -129 565 -29 603
rect 29 637 129 675
rect 29 603 45 637
rect 113 603 129 637
rect 29 565 129 603
rect 187 637 287 675
rect 187 603 203 637
rect 271 603 287 637
rect 187 565 287 603
rect 345 637 445 675
rect 345 603 361 637
rect 429 603 445 637
rect 345 565 445 603
rect 503 637 603 675
rect 503 603 519 637
rect 587 603 603 637
rect 503 565 603 603
rect 661 637 761 675
rect 661 603 677 637
rect 745 603 761 637
rect 661 565 761 603
rect 819 637 919 675
rect 819 603 835 637
rect 903 603 919 637
rect 819 565 919 603
rect 977 637 1077 675
rect 977 603 993 637
rect 1061 603 1077 637
rect 977 565 1077 603
rect 1135 637 1235 675
rect 1135 603 1151 637
rect 1219 603 1235 637
rect 1135 565 1235 603
rect 1293 637 1393 675
rect 1293 603 1309 637
rect 1377 603 1393 637
rect 1293 565 1393 603
rect 1451 637 1551 675
rect 1451 603 1467 637
rect 1535 603 1551 637
rect 1451 565 1551 603
rect -1551 327 -1451 365
rect -1551 293 -1535 327
rect -1467 293 -1451 327
rect -1551 255 -1451 293
rect -1393 327 -1293 365
rect -1393 293 -1377 327
rect -1309 293 -1293 327
rect -1393 255 -1293 293
rect -1235 327 -1135 365
rect -1235 293 -1219 327
rect -1151 293 -1135 327
rect -1235 255 -1135 293
rect -1077 327 -977 365
rect -1077 293 -1061 327
rect -993 293 -977 327
rect -1077 255 -977 293
rect -919 327 -819 365
rect -919 293 -903 327
rect -835 293 -819 327
rect -919 255 -819 293
rect -761 327 -661 365
rect -761 293 -745 327
rect -677 293 -661 327
rect -761 255 -661 293
rect -603 327 -503 365
rect -603 293 -587 327
rect -519 293 -503 327
rect -603 255 -503 293
rect -445 327 -345 365
rect -445 293 -429 327
rect -361 293 -345 327
rect -445 255 -345 293
rect -287 327 -187 365
rect -287 293 -271 327
rect -203 293 -187 327
rect -287 255 -187 293
rect -129 327 -29 365
rect -129 293 -113 327
rect -45 293 -29 327
rect -129 255 -29 293
rect 29 327 129 365
rect 29 293 45 327
rect 113 293 129 327
rect 29 255 129 293
rect 187 327 287 365
rect 187 293 203 327
rect 271 293 287 327
rect 187 255 287 293
rect 345 327 445 365
rect 345 293 361 327
rect 429 293 445 327
rect 345 255 445 293
rect 503 327 603 365
rect 503 293 519 327
rect 587 293 603 327
rect 503 255 603 293
rect 661 327 761 365
rect 661 293 677 327
rect 745 293 761 327
rect 661 255 761 293
rect 819 327 919 365
rect 819 293 835 327
rect 903 293 919 327
rect 819 255 919 293
rect 977 327 1077 365
rect 977 293 993 327
rect 1061 293 1077 327
rect 977 255 1077 293
rect 1135 327 1235 365
rect 1135 293 1151 327
rect 1219 293 1235 327
rect 1135 255 1235 293
rect 1293 327 1393 365
rect 1293 293 1309 327
rect 1377 293 1393 327
rect 1293 255 1393 293
rect 1451 327 1551 365
rect 1451 293 1467 327
rect 1535 293 1551 327
rect 1451 255 1551 293
rect -1551 17 -1451 55
rect -1551 -17 -1535 17
rect -1467 -17 -1451 17
rect -1551 -55 -1451 -17
rect -1393 17 -1293 55
rect -1393 -17 -1377 17
rect -1309 -17 -1293 17
rect -1393 -55 -1293 -17
rect -1235 17 -1135 55
rect -1235 -17 -1219 17
rect -1151 -17 -1135 17
rect -1235 -55 -1135 -17
rect -1077 17 -977 55
rect -1077 -17 -1061 17
rect -993 -17 -977 17
rect -1077 -55 -977 -17
rect -919 17 -819 55
rect -919 -17 -903 17
rect -835 -17 -819 17
rect -919 -55 -819 -17
rect -761 17 -661 55
rect -761 -17 -745 17
rect -677 -17 -661 17
rect -761 -55 -661 -17
rect -603 17 -503 55
rect -603 -17 -587 17
rect -519 -17 -503 17
rect -603 -55 -503 -17
rect -445 17 -345 55
rect -445 -17 -429 17
rect -361 -17 -345 17
rect -445 -55 -345 -17
rect -287 17 -187 55
rect -287 -17 -271 17
rect -203 -17 -187 17
rect -287 -55 -187 -17
rect -129 17 -29 55
rect -129 -17 -113 17
rect -45 -17 -29 17
rect -129 -55 -29 -17
rect 29 17 129 55
rect 29 -17 45 17
rect 113 -17 129 17
rect 29 -55 129 -17
rect 187 17 287 55
rect 187 -17 203 17
rect 271 -17 287 17
rect 187 -55 287 -17
rect 345 17 445 55
rect 345 -17 361 17
rect 429 -17 445 17
rect 345 -55 445 -17
rect 503 17 603 55
rect 503 -17 519 17
rect 587 -17 603 17
rect 503 -55 603 -17
rect 661 17 761 55
rect 661 -17 677 17
rect 745 -17 761 17
rect 661 -55 761 -17
rect 819 17 919 55
rect 819 -17 835 17
rect 903 -17 919 17
rect 819 -55 919 -17
rect 977 17 1077 55
rect 977 -17 993 17
rect 1061 -17 1077 17
rect 977 -55 1077 -17
rect 1135 17 1235 55
rect 1135 -17 1151 17
rect 1219 -17 1235 17
rect 1135 -55 1235 -17
rect 1293 17 1393 55
rect 1293 -17 1309 17
rect 1377 -17 1393 17
rect 1293 -55 1393 -17
rect 1451 17 1551 55
rect 1451 -17 1467 17
rect 1535 -17 1551 17
rect 1451 -55 1551 -17
rect -1551 -293 -1451 -255
rect -1551 -327 -1535 -293
rect -1467 -327 -1451 -293
rect -1551 -365 -1451 -327
rect -1393 -293 -1293 -255
rect -1393 -327 -1377 -293
rect -1309 -327 -1293 -293
rect -1393 -365 -1293 -327
rect -1235 -293 -1135 -255
rect -1235 -327 -1219 -293
rect -1151 -327 -1135 -293
rect -1235 -365 -1135 -327
rect -1077 -293 -977 -255
rect -1077 -327 -1061 -293
rect -993 -327 -977 -293
rect -1077 -365 -977 -327
rect -919 -293 -819 -255
rect -919 -327 -903 -293
rect -835 -327 -819 -293
rect -919 -365 -819 -327
rect -761 -293 -661 -255
rect -761 -327 -745 -293
rect -677 -327 -661 -293
rect -761 -365 -661 -327
rect -603 -293 -503 -255
rect -603 -327 -587 -293
rect -519 -327 -503 -293
rect -603 -365 -503 -327
rect -445 -293 -345 -255
rect -445 -327 -429 -293
rect -361 -327 -345 -293
rect -445 -365 -345 -327
rect -287 -293 -187 -255
rect -287 -327 -271 -293
rect -203 -327 -187 -293
rect -287 -365 -187 -327
rect -129 -293 -29 -255
rect -129 -327 -113 -293
rect -45 -327 -29 -293
rect -129 -365 -29 -327
rect 29 -293 129 -255
rect 29 -327 45 -293
rect 113 -327 129 -293
rect 29 -365 129 -327
rect 187 -293 287 -255
rect 187 -327 203 -293
rect 271 -327 287 -293
rect 187 -365 287 -327
rect 345 -293 445 -255
rect 345 -327 361 -293
rect 429 -327 445 -293
rect 345 -365 445 -327
rect 503 -293 603 -255
rect 503 -327 519 -293
rect 587 -327 603 -293
rect 503 -365 603 -327
rect 661 -293 761 -255
rect 661 -327 677 -293
rect 745 -327 761 -293
rect 661 -365 761 -327
rect 819 -293 919 -255
rect 819 -327 835 -293
rect 903 -327 919 -293
rect 819 -365 919 -327
rect 977 -293 1077 -255
rect 977 -327 993 -293
rect 1061 -327 1077 -293
rect 977 -365 1077 -327
rect 1135 -293 1235 -255
rect 1135 -327 1151 -293
rect 1219 -327 1235 -293
rect 1135 -365 1235 -327
rect 1293 -293 1393 -255
rect 1293 -327 1309 -293
rect 1377 -327 1393 -293
rect 1293 -365 1393 -327
rect 1451 -293 1551 -255
rect 1451 -327 1467 -293
rect 1535 -327 1551 -293
rect 1451 -365 1551 -327
rect -1551 -603 -1451 -565
rect -1551 -637 -1535 -603
rect -1467 -637 -1451 -603
rect -1551 -675 -1451 -637
rect -1393 -603 -1293 -565
rect -1393 -637 -1377 -603
rect -1309 -637 -1293 -603
rect -1393 -675 -1293 -637
rect -1235 -603 -1135 -565
rect -1235 -637 -1219 -603
rect -1151 -637 -1135 -603
rect -1235 -675 -1135 -637
rect -1077 -603 -977 -565
rect -1077 -637 -1061 -603
rect -993 -637 -977 -603
rect -1077 -675 -977 -637
rect -919 -603 -819 -565
rect -919 -637 -903 -603
rect -835 -637 -819 -603
rect -919 -675 -819 -637
rect -761 -603 -661 -565
rect -761 -637 -745 -603
rect -677 -637 -661 -603
rect -761 -675 -661 -637
rect -603 -603 -503 -565
rect -603 -637 -587 -603
rect -519 -637 -503 -603
rect -603 -675 -503 -637
rect -445 -603 -345 -565
rect -445 -637 -429 -603
rect -361 -637 -345 -603
rect -445 -675 -345 -637
rect -287 -603 -187 -565
rect -287 -637 -271 -603
rect -203 -637 -187 -603
rect -287 -675 -187 -637
rect -129 -603 -29 -565
rect -129 -637 -113 -603
rect -45 -637 -29 -603
rect -129 -675 -29 -637
rect 29 -603 129 -565
rect 29 -637 45 -603
rect 113 -637 129 -603
rect 29 -675 129 -637
rect 187 -603 287 -565
rect 187 -637 203 -603
rect 271 -637 287 -603
rect 187 -675 287 -637
rect 345 -603 445 -565
rect 345 -637 361 -603
rect 429 -637 445 -603
rect 345 -675 445 -637
rect 503 -603 603 -565
rect 503 -637 519 -603
rect 587 -637 603 -603
rect 503 -675 603 -637
rect 661 -603 761 -565
rect 661 -637 677 -603
rect 745 -637 761 -603
rect 661 -675 761 -637
rect 819 -603 919 -565
rect 819 -637 835 -603
rect 903 -637 919 -603
rect 819 -675 919 -637
rect 977 -603 1077 -565
rect 977 -637 993 -603
rect 1061 -637 1077 -603
rect 977 -675 1077 -637
rect 1135 -603 1235 -565
rect 1135 -637 1151 -603
rect 1219 -637 1235 -603
rect 1135 -675 1235 -637
rect 1293 -603 1393 -565
rect 1293 -637 1309 -603
rect 1377 -637 1393 -603
rect 1293 -675 1393 -637
rect 1451 -603 1551 -565
rect 1451 -637 1467 -603
rect 1535 -637 1551 -603
rect 1451 -675 1551 -637
rect -1551 -913 -1451 -875
rect -1551 -947 -1535 -913
rect -1467 -947 -1451 -913
rect -1551 -985 -1451 -947
rect -1393 -913 -1293 -875
rect -1393 -947 -1377 -913
rect -1309 -947 -1293 -913
rect -1393 -985 -1293 -947
rect -1235 -913 -1135 -875
rect -1235 -947 -1219 -913
rect -1151 -947 -1135 -913
rect -1235 -985 -1135 -947
rect -1077 -913 -977 -875
rect -1077 -947 -1061 -913
rect -993 -947 -977 -913
rect -1077 -985 -977 -947
rect -919 -913 -819 -875
rect -919 -947 -903 -913
rect -835 -947 -819 -913
rect -919 -985 -819 -947
rect -761 -913 -661 -875
rect -761 -947 -745 -913
rect -677 -947 -661 -913
rect -761 -985 -661 -947
rect -603 -913 -503 -875
rect -603 -947 -587 -913
rect -519 -947 -503 -913
rect -603 -985 -503 -947
rect -445 -913 -345 -875
rect -445 -947 -429 -913
rect -361 -947 -345 -913
rect -445 -985 -345 -947
rect -287 -913 -187 -875
rect -287 -947 -271 -913
rect -203 -947 -187 -913
rect -287 -985 -187 -947
rect -129 -913 -29 -875
rect -129 -947 -113 -913
rect -45 -947 -29 -913
rect -129 -985 -29 -947
rect 29 -913 129 -875
rect 29 -947 45 -913
rect 113 -947 129 -913
rect 29 -985 129 -947
rect 187 -913 287 -875
rect 187 -947 203 -913
rect 271 -947 287 -913
rect 187 -985 287 -947
rect 345 -913 445 -875
rect 345 -947 361 -913
rect 429 -947 445 -913
rect 345 -985 445 -947
rect 503 -913 603 -875
rect 503 -947 519 -913
rect 587 -947 603 -913
rect 503 -985 603 -947
rect 661 -913 761 -875
rect 661 -947 677 -913
rect 745 -947 761 -913
rect 661 -985 761 -947
rect 819 -913 919 -875
rect 819 -947 835 -913
rect 903 -947 919 -913
rect 819 -985 919 -947
rect 977 -913 1077 -875
rect 977 -947 993 -913
rect 1061 -947 1077 -913
rect 977 -985 1077 -947
rect 1135 -913 1235 -875
rect 1135 -947 1151 -913
rect 1219 -947 1235 -913
rect 1135 -985 1235 -947
rect 1293 -913 1393 -875
rect 1293 -947 1309 -913
rect 1377 -947 1393 -913
rect 1293 -985 1393 -947
rect 1451 -913 1551 -875
rect 1451 -947 1467 -913
rect 1535 -947 1551 -913
rect 1451 -985 1551 -947
rect -1551 -1223 -1451 -1185
rect -1551 -1257 -1535 -1223
rect -1467 -1257 -1451 -1223
rect -1551 -1295 -1451 -1257
rect -1393 -1223 -1293 -1185
rect -1393 -1257 -1377 -1223
rect -1309 -1257 -1293 -1223
rect -1393 -1295 -1293 -1257
rect -1235 -1223 -1135 -1185
rect -1235 -1257 -1219 -1223
rect -1151 -1257 -1135 -1223
rect -1235 -1295 -1135 -1257
rect -1077 -1223 -977 -1185
rect -1077 -1257 -1061 -1223
rect -993 -1257 -977 -1223
rect -1077 -1295 -977 -1257
rect -919 -1223 -819 -1185
rect -919 -1257 -903 -1223
rect -835 -1257 -819 -1223
rect -919 -1295 -819 -1257
rect -761 -1223 -661 -1185
rect -761 -1257 -745 -1223
rect -677 -1257 -661 -1223
rect -761 -1295 -661 -1257
rect -603 -1223 -503 -1185
rect -603 -1257 -587 -1223
rect -519 -1257 -503 -1223
rect -603 -1295 -503 -1257
rect -445 -1223 -345 -1185
rect -445 -1257 -429 -1223
rect -361 -1257 -345 -1223
rect -445 -1295 -345 -1257
rect -287 -1223 -187 -1185
rect -287 -1257 -271 -1223
rect -203 -1257 -187 -1223
rect -287 -1295 -187 -1257
rect -129 -1223 -29 -1185
rect -129 -1257 -113 -1223
rect -45 -1257 -29 -1223
rect -129 -1295 -29 -1257
rect 29 -1223 129 -1185
rect 29 -1257 45 -1223
rect 113 -1257 129 -1223
rect 29 -1295 129 -1257
rect 187 -1223 287 -1185
rect 187 -1257 203 -1223
rect 271 -1257 287 -1223
rect 187 -1295 287 -1257
rect 345 -1223 445 -1185
rect 345 -1257 361 -1223
rect 429 -1257 445 -1223
rect 345 -1295 445 -1257
rect 503 -1223 603 -1185
rect 503 -1257 519 -1223
rect 587 -1257 603 -1223
rect 503 -1295 603 -1257
rect 661 -1223 761 -1185
rect 661 -1257 677 -1223
rect 745 -1257 761 -1223
rect 661 -1295 761 -1257
rect 819 -1223 919 -1185
rect 819 -1257 835 -1223
rect 903 -1257 919 -1223
rect 819 -1295 919 -1257
rect 977 -1223 1077 -1185
rect 977 -1257 993 -1223
rect 1061 -1257 1077 -1223
rect 977 -1295 1077 -1257
rect 1135 -1223 1235 -1185
rect 1135 -1257 1151 -1223
rect 1219 -1257 1235 -1223
rect 1135 -1295 1235 -1257
rect 1293 -1223 1393 -1185
rect 1293 -1257 1309 -1223
rect 1377 -1257 1393 -1223
rect 1293 -1295 1393 -1257
rect 1451 -1223 1551 -1185
rect 1451 -1257 1467 -1223
rect 1535 -1257 1551 -1223
rect 1451 -1295 1551 -1257
rect -1551 -1533 -1451 -1495
rect -1551 -1567 -1535 -1533
rect -1467 -1567 -1451 -1533
rect -1551 -1583 -1451 -1567
rect -1393 -1533 -1293 -1495
rect -1393 -1567 -1377 -1533
rect -1309 -1567 -1293 -1533
rect -1393 -1583 -1293 -1567
rect -1235 -1533 -1135 -1495
rect -1235 -1567 -1219 -1533
rect -1151 -1567 -1135 -1533
rect -1235 -1583 -1135 -1567
rect -1077 -1533 -977 -1495
rect -1077 -1567 -1061 -1533
rect -993 -1567 -977 -1533
rect -1077 -1583 -977 -1567
rect -919 -1533 -819 -1495
rect -919 -1567 -903 -1533
rect -835 -1567 -819 -1533
rect -919 -1583 -819 -1567
rect -761 -1533 -661 -1495
rect -761 -1567 -745 -1533
rect -677 -1567 -661 -1533
rect -761 -1583 -661 -1567
rect -603 -1533 -503 -1495
rect -603 -1567 -587 -1533
rect -519 -1567 -503 -1533
rect -603 -1583 -503 -1567
rect -445 -1533 -345 -1495
rect -445 -1567 -429 -1533
rect -361 -1567 -345 -1533
rect -445 -1583 -345 -1567
rect -287 -1533 -187 -1495
rect -287 -1567 -271 -1533
rect -203 -1567 -187 -1533
rect -287 -1583 -187 -1567
rect -129 -1533 -29 -1495
rect -129 -1567 -113 -1533
rect -45 -1567 -29 -1533
rect -129 -1583 -29 -1567
rect 29 -1533 129 -1495
rect 29 -1567 45 -1533
rect 113 -1567 129 -1533
rect 29 -1583 129 -1567
rect 187 -1533 287 -1495
rect 187 -1567 203 -1533
rect 271 -1567 287 -1533
rect 187 -1583 287 -1567
rect 345 -1533 445 -1495
rect 345 -1567 361 -1533
rect 429 -1567 445 -1533
rect 345 -1583 445 -1567
rect 503 -1533 603 -1495
rect 503 -1567 519 -1533
rect 587 -1567 603 -1533
rect 503 -1583 603 -1567
rect 661 -1533 761 -1495
rect 661 -1567 677 -1533
rect 745 -1567 761 -1533
rect 661 -1583 761 -1567
rect 819 -1533 919 -1495
rect 819 -1567 835 -1533
rect 903 -1567 919 -1533
rect 819 -1583 919 -1567
rect 977 -1533 1077 -1495
rect 977 -1567 993 -1533
rect 1061 -1567 1077 -1533
rect 977 -1583 1077 -1567
rect 1135 -1533 1235 -1495
rect 1135 -1567 1151 -1533
rect 1219 -1567 1235 -1533
rect 1135 -1583 1235 -1567
rect 1293 -1533 1393 -1495
rect 1293 -1567 1309 -1533
rect 1377 -1567 1393 -1533
rect 1293 -1583 1393 -1567
rect 1451 -1533 1551 -1495
rect 1451 -1567 1467 -1533
rect 1535 -1567 1551 -1533
rect 1451 -1583 1551 -1567
<< polycont >>
rect -1535 1533 -1467 1567
rect -1377 1533 -1309 1567
rect -1219 1533 -1151 1567
rect -1061 1533 -993 1567
rect -903 1533 -835 1567
rect -745 1533 -677 1567
rect -587 1533 -519 1567
rect -429 1533 -361 1567
rect -271 1533 -203 1567
rect -113 1533 -45 1567
rect 45 1533 113 1567
rect 203 1533 271 1567
rect 361 1533 429 1567
rect 519 1533 587 1567
rect 677 1533 745 1567
rect 835 1533 903 1567
rect 993 1533 1061 1567
rect 1151 1533 1219 1567
rect 1309 1533 1377 1567
rect 1467 1533 1535 1567
rect -1535 1223 -1467 1257
rect -1377 1223 -1309 1257
rect -1219 1223 -1151 1257
rect -1061 1223 -993 1257
rect -903 1223 -835 1257
rect -745 1223 -677 1257
rect -587 1223 -519 1257
rect -429 1223 -361 1257
rect -271 1223 -203 1257
rect -113 1223 -45 1257
rect 45 1223 113 1257
rect 203 1223 271 1257
rect 361 1223 429 1257
rect 519 1223 587 1257
rect 677 1223 745 1257
rect 835 1223 903 1257
rect 993 1223 1061 1257
rect 1151 1223 1219 1257
rect 1309 1223 1377 1257
rect 1467 1223 1535 1257
rect -1535 913 -1467 947
rect -1377 913 -1309 947
rect -1219 913 -1151 947
rect -1061 913 -993 947
rect -903 913 -835 947
rect -745 913 -677 947
rect -587 913 -519 947
rect -429 913 -361 947
rect -271 913 -203 947
rect -113 913 -45 947
rect 45 913 113 947
rect 203 913 271 947
rect 361 913 429 947
rect 519 913 587 947
rect 677 913 745 947
rect 835 913 903 947
rect 993 913 1061 947
rect 1151 913 1219 947
rect 1309 913 1377 947
rect 1467 913 1535 947
rect -1535 603 -1467 637
rect -1377 603 -1309 637
rect -1219 603 -1151 637
rect -1061 603 -993 637
rect -903 603 -835 637
rect -745 603 -677 637
rect -587 603 -519 637
rect -429 603 -361 637
rect -271 603 -203 637
rect -113 603 -45 637
rect 45 603 113 637
rect 203 603 271 637
rect 361 603 429 637
rect 519 603 587 637
rect 677 603 745 637
rect 835 603 903 637
rect 993 603 1061 637
rect 1151 603 1219 637
rect 1309 603 1377 637
rect 1467 603 1535 637
rect -1535 293 -1467 327
rect -1377 293 -1309 327
rect -1219 293 -1151 327
rect -1061 293 -993 327
rect -903 293 -835 327
rect -745 293 -677 327
rect -587 293 -519 327
rect -429 293 -361 327
rect -271 293 -203 327
rect -113 293 -45 327
rect 45 293 113 327
rect 203 293 271 327
rect 361 293 429 327
rect 519 293 587 327
rect 677 293 745 327
rect 835 293 903 327
rect 993 293 1061 327
rect 1151 293 1219 327
rect 1309 293 1377 327
rect 1467 293 1535 327
rect -1535 -17 -1467 17
rect -1377 -17 -1309 17
rect -1219 -17 -1151 17
rect -1061 -17 -993 17
rect -903 -17 -835 17
rect -745 -17 -677 17
rect -587 -17 -519 17
rect -429 -17 -361 17
rect -271 -17 -203 17
rect -113 -17 -45 17
rect 45 -17 113 17
rect 203 -17 271 17
rect 361 -17 429 17
rect 519 -17 587 17
rect 677 -17 745 17
rect 835 -17 903 17
rect 993 -17 1061 17
rect 1151 -17 1219 17
rect 1309 -17 1377 17
rect 1467 -17 1535 17
rect -1535 -327 -1467 -293
rect -1377 -327 -1309 -293
rect -1219 -327 -1151 -293
rect -1061 -327 -993 -293
rect -903 -327 -835 -293
rect -745 -327 -677 -293
rect -587 -327 -519 -293
rect -429 -327 -361 -293
rect -271 -327 -203 -293
rect -113 -327 -45 -293
rect 45 -327 113 -293
rect 203 -327 271 -293
rect 361 -327 429 -293
rect 519 -327 587 -293
rect 677 -327 745 -293
rect 835 -327 903 -293
rect 993 -327 1061 -293
rect 1151 -327 1219 -293
rect 1309 -327 1377 -293
rect 1467 -327 1535 -293
rect -1535 -637 -1467 -603
rect -1377 -637 -1309 -603
rect -1219 -637 -1151 -603
rect -1061 -637 -993 -603
rect -903 -637 -835 -603
rect -745 -637 -677 -603
rect -587 -637 -519 -603
rect -429 -637 -361 -603
rect -271 -637 -203 -603
rect -113 -637 -45 -603
rect 45 -637 113 -603
rect 203 -637 271 -603
rect 361 -637 429 -603
rect 519 -637 587 -603
rect 677 -637 745 -603
rect 835 -637 903 -603
rect 993 -637 1061 -603
rect 1151 -637 1219 -603
rect 1309 -637 1377 -603
rect 1467 -637 1535 -603
rect -1535 -947 -1467 -913
rect -1377 -947 -1309 -913
rect -1219 -947 -1151 -913
rect -1061 -947 -993 -913
rect -903 -947 -835 -913
rect -745 -947 -677 -913
rect -587 -947 -519 -913
rect -429 -947 -361 -913
rect -271 -947 -203 -913
rect -113 -947 -45 -913
rect 45 -947 113 -913
rect 203 -947 271 -913
rect 361 -947 429 -913
rect 519 -947 587 -913
rect 677 -947 745 -913
rect 835 -947 903 -913
rect 993 -947 1061 -913
rect 1151 -947 1219 -913
rect 1309 -947 1377 -913
rect 1467 -947 1535 -913
rect -1535 -1257 -1467 -1223
rect -1377 -1257 -1309 -1223
rect -1219 -1257 -1151 -1223
rect -1061 -1257 -993 -1223
rect -903 -1257 -835 -1223
rect -745 -1257 -677 -1223
rect -587 -1257 -519 -1223
rect -429 -1257 -361 -1223
rect -271 -1257 -203 -1223
rect -113 -1257 -45 -1223
rect 45 -1257 113 -1223
rect 203 -1257 271 -1223
rect 361 -1257 429 -1223
rect 519 -1257 587 -1223
rect 677 -1257 745 -1223
rect 835 -1257 903 -1223
rect 993 -1257 1061 -1223
rect 1151 -1257 1219 -1223
rect 1309 -1257 1377 -1223
rect 1467 -1257 1535 -1223
rect -1535 -1567 -1467 -1533
rect -1377 -1567 -1309 -1533
rect -1219 -1567 -1151 -1533
rect -1061 -1567 -993 -1533
rect -903 -1567 -835 -1533
rect -745 -1567 -677 -1533
rect -587 -1567 -519 -1533
rect -429 -1567 -361 -1533
rect -271 -1567 -203 -1533
rect -113 -1567 -45 -1533
rect 45 -1567 113 -1533
rect 203 -1567 271 -1533
rect 361 -1567 429 -1533
rect 519 -1567 587 -1533
rect 677 -1567 745 -1533
rect 835 -1567 903 -1533
rect 993 -1567 1061 -1533
rect 1151 -1567 1219 -1533
rect 1309 -1567 1377 -1533
rect 1467 -1567 1535 -1533
<< locali >>
rect -1731 1671 -1635 1705
rect 1635 1671 1731 1705
rect -1731 1609 -1697 1671
rect 1697 1609 1731 1671
rect -1551 1533 -1535 1567
rect -1467 1533 -1451 1567
rect -1393 1533 -1377 1567
rect -1309 1533 -1293 1567
rect -1235 1533 -1219 1567
rect -1151 1533 -1135 1567
rect -1077 1533 -1061 1567
rect -993 1533 -977 1567
rect -919 1533 -903 1567
rect -835 1533 -819 1567
rect -761 1533 -745 1567
rect -677 1533 -661 1567
rect -603 1533 -587 1567
rect -519 1533 -503 1567
rect -445 1533 -429 1567
rect -361 1533 -345 1567
rect -287 1533 -271 1567
rect -203 1533 -187 1567
rect -129 1533 -113 1567
rect -45 1533 -29 1567
rect 29 1533 45 1567
rect 113 1533 129 1567
rect 187 1533 203 1567
rect 271 1533 287 1567
rect 345 1533 361 1567
rect 429 1533 445 1567
rect 503 1533 519 1567
rect 587 1533 603 1567
rect 661 1533 677 1567
rect 745 1533 761 1567
rect 819 1533 835 1567
rect 903 1533 919 1567
rect 977 1533 993 1567
rect 1061 1533 1077 1567
rect 1135 1533 1151 1567
rect 1219 1533 1235 1567
rect 1293 1533 1309 1567
rect 1377 1533 1393 1567
rect 1451 1533 1467 1567
rect 1535 1533 1551 1567
rect -1597 1483 -1563 1499
rect -1597 1291 -1563 1307
rect -1439 1483 -1405 1499
rect -1439 1291 -1405 1307
rect -1281 1483 -1247 1499
rect -1281 1291 -1247 1307
rect -1123 1483 -1089 1499
rect -1123 1291 -1089 1307
rect -965 1483 -931 1499
rect -965 1291 -931 1307
rect -807 1483 -773 1499
rect -807 1291 -773 1307
rect -649 1483 -615 1499
rect -649 1291 -615 1307
rect -491 1483 -457 1499
rect -491 1291 -457 1307
rect -333 1483 -299 1499
rect -333 1291 -299 1307
rect -175 1483 -141 1499
rect -175 1291 -141 1307
rect -17 1483 17 1499
rect -17 1291 17 1307
rect 141 1483 175 1499
rect 141 1291 175 1307
rect 299 1483 333 1499
rect 299 1291 333 1307
rect 457 1483 491 1499
rect 457 1291 491 1307
rect 615 1483 649 1499
rect 615 1291 649 1307
rect 773 1483 807 1499
rect 773 1291 807 1307
rect 931 1483 965 1499
rect 931 1291 965 1307
rect 1089 1483 1123 1499
rect 1089 1291 1123 1307
rect 1247 1483 1281 1499
rect 1247 1291 1281 1307
rect 1405 1483 1439 1499
rect 1405 1291 1439 1307
rect 1563 1483 1597 1499
rect 1563 1291 1597 1307
rect -1551 1223 -1535 1257
rect -1467 1223 -1451 1257
rect -1393 1223 -1377 1257
rect -1309 1223 -1293 1257
rect -1235 1223 -1219 1257
rect -1151 1223 -1135 1257
rect -1077 1223 -1061 1257
rect -993 1223 -977 1257
rect -919 1223 -903 1257
rect -835 1223 -819 1257
rect -761 1223 -745 1257
rect -677 1223 -661 1257
rect -603 1223 -587 1257
rect -519 1223 -503 1257
rect -445 1223 -429 1257
rect -361 1223 -345 1257
rect -287 1223 -271 1257
rect -203 1223 -187 1257
rect -129 1223 -113 1257
rect -45 1223 -29 1257
rect 29 1223 45 1257
rect 113 1223 129 1257
rect 187 1223 203 1257
rect 271 1223 287 1257
rect 345 1223 361 1257
rect 429 1223 445 1257
rect 503 1223 519 1257
rect 587 1223 603 1257
rect 661 1223 677 1257
rect 745 1223 761 1257
rect 819 1223 835 1257
rect 903 1223 919 1257
rect 977 1223 993 1257
rect 1061 1223 1077 1257
rect 1135 1223 1151 1257
rect 1219 1223 1235 1257
rect 1293 1223 1309 1257
rect 1377 1223 1393 1257
rect 1451 1223 1467 1257
rect 1535 1223 1551 1257
rect -1597 1173 -1563 1189
rect -1597 981 -1563 997
rect -1439 1173 -1405 1189
rect -1439 981 -1405 997
rect -1281 1173 -1247 1189
rect -1281 981 -1247 997
rect -1123 1173 -1089 1189
rect -1123 981 -1089 997
rect -965 1173 -931 1189
rect -965 981 -931 997
rect -807 1173 -773 1189
rect -807 981 -773 997
rect -649 1173 -615 1189
rect -649 981 -615 997
rect -491 1173 -457 1189
rect -491 981 -457 997
rect -333 1173 -299 1189
rect -333 981 -299 997
rect -175 1173 -141 1189
rect -175 981 -141 997
rect -17 1173 17 1189
rect -17 981 17 997
rect 141 1173 175 1189
rect 141 981 175 997
rect 299 1173 333 1189
rect 299 981 333 997
rect 457 1173 491 1189
rect 457 981 491 997
rect 615 1173 649 1189
rect 615 981 649 997
rect 773 1173 807 1189
rect 773 981 807 997
rect 931 1173 965 1189
rect 931 981 965 997
rect 1089 1173 1123 1189
rect 1089 981 1123 997
rect 1247 1173 1281 1189
rect 1247 981 1281 997
rect 1405 1173 1439 1189
rect 1405 981 1439 997
rect 1563 1173 1597 1189
rect 1563 981 1597 997
rect -1551 913 -1535 947
rect -1467 913 -1451 947
rect -1393 913 -1377 947
rect -1309 913 -1293 947
rect -1235 913 -1219 947
rect -1151 913 -1135 947
rect -1077 913 -1061 947
rect -993 913 -977 947
rect -919 913 -903 947
rect -835 913 -819 947
rect -761 913 -745 947
rect -677 913 -661 947
rect -603 913 -587 947
rect -519 913 -503 947
rect -445 913 -429 947
rect -361 913 -345 947
rect -287 913 -271 947
rect -203 913 -187 947
rect -129 913 -113 947
rect -45 913 -29 947
rect 29 913 45 947
rect 113 913 129 947
rect 187 913 203 947
rect 271 913 287 947
rect 345 913 361 947
rect 429 913 445 947
rect 503 913 519 947
rect 587 913 603 947
rect 661 913 677 947
rect 745 913 761 947
rect 819 913 835 947
rect 903 913 919 947
rect 977 913 993 947
rect 1061 913 1077 947
rect 1135 913 1151 947
rect 1219 913 1235 947
rect 1293 913 1309 947
rect 1377 913 1393 947
rect 1451 913 1467 947
rect 1535 913 1551 947
rect -1597 863 -1563 879
rect -1597 671 -1563 687
rect -1439 863 -1405 879
rect -1439 671 -1405 687
rect -1281 863 -1247 879
rect -1281 671 -1247 687
rect -1123 863 -1089 879
rect -1123 671 -1089 687
rect -965 863 -931 879
rect -965 671 -931 687
rect -807 863 -773 879
rect -807 671 -773 687
rect -649 863 -615 879
rect -649 671 -615 687
rect -491 863 -457 879
rect -491 671 -457 687
rect -333 863 -299 879
rect -333 671 -299 687
rect -175 863 -141 879
rect -175 671 -141 687
rect -17 863 17 879
rect -17 671 17 687
rect 141 863 175 879
rect 141 671 175 687
rect 299 863 333 879
rect 299 671 333 687
rect 457 863 491 879
rect 457 671 491 687
rect 615 863 649 879
rect 615 671 649 687
rect 773 863 807 879
rect 773 671 807 687
rect 931 863 965 879
rect 931 671 965 687
rect 1089 863 1123 879
rect 1089 671 1123 687
rect 1247 863 1281 879
rect 1247 671 1281 687
rect 1405 863 1439 879
rect 1405 671 1439 687
rect 1563 863 1597 879
rect 1563 671 1597 687
rect -1551 603 -1535 637
rect -1467 603 -1451 637
rect -1393 603 -1377 637
rect -1309 603 -1293 637
rect -1235 603 -1219 637
rect -1151 603 -1135 637
rect -1077 603 -1061 637
rect -993 603 -977 637
rect -919 603 -903 637
rect -835 603 -819 637
rect -761 603 -745 637
rect -677 603 -661 637
rect -603 603 -587 637
rect -519 603 -503 637
rect -445 603 -429 637
rect -361 603 -345 637
rect -287 603 -271 637
rect -203 603 -187 637
rect -129 603 -113 637
rect -45 603 -29 637
rect 29 603 45 637
rect 113 603 129 637
rect 187 603 203 637
rect 271 603 287 637
rect 345 603 361 637
rect 429 603 445 637
rect 503 603 519 637
rect 587 603 603 637
rect 661 603 677 637
rect 745 603 761 637
rect 819 603 835 637
rect 903 603 919 637
rect 977 603 993 637
rect 1061 603 1077 637
rect 1135 603 1151 637
rect 1219 603 1235 637
rect 1293 603 1309 637
rect 1377 603 1393 637
rect 1451 603 1467 637
rect 1535 603 1551 637
rect -1597 553 -1563 569
rect -1597 361 -1563 377
rect -1439 553 -1405 569
rect -1439 361 -1405 377
rect -1281 553 -1247 569
rect -1281 361 -1247 377
rect -1123 553 -1089 569
rect -1123 361 -1089 377
rect -965 553 -931 569
rect -965 361 -931 377
rect -807 553 -773 569
rect -807 361 -773 377
rect -649 553 -615 569
rect -649 361 -615 377
rect -491 553 -457 569
rect -491 361 -457 377
rect -333 553 -299 569
rect -333 361 -299 377
rect -175 553 -141 569
rect -175 361 -141 377
rect -17 553 17 569
rect -17 361 17 377
rect 141 553 175 569
rect 141 361 175 377
rect 299 553 333 569
rect 299 361 333 377
rect 457 553 491 569
rect 457 361 491 377
rect 615 553 649 569
rect 615 361 649 377
rect 773 553 807 569
rect 773 361 807 377
rect 931 553 965 569
rect 931 361 965 377
rect 1089 553 1123 569
rect 1089 361 1123 377
rect 1247 553 1281 569
rect 1247 361 1281 377
rect 1405 553 1439 569
rect 1405 361 1439 377
rect 1563 553 1597 569
rect 1563 361 1597 377
rect -1551 293 -1535 327
rect -1467 293 -1451 327
rect -1393 293 -1377 327
rect -1309 293 -1293 327
rect -1235 293 -1219 327
rect -1151 293 -1135 327
rect -1077 293 -1061 327
rect -993 293 -977 327
rect -919 293 -903 327
rect -835 293 -819 327
rect -761 293 -745 327
rect -677 293 -661 327
rect -603 293 -587 327
rect -519 293 -503 327
rect -445 293 -429 327
rect -361 293 -345 327
rect -287 293 -271 327
rect -203 293 -187 327
rect -129 293 -113 327
rect -45 293 -29 327
rect 29 293 45 327
rect 113 293 129 327
rect 187 293 203 327
rect 271 293 287 327
rect 345 293 361 327
rect 429 293 445 327
rect 503 293 519 327
rect 587 293 603 327
rect 661 293 677 327
rect 745 293 761 327
rect 819 293 835 327
rect 903 293 919 327
rect 977 293 993 327
rect 1061 293 1077 327
rect 1135 293 1151 327
rect 1219 293 1235 327
rect 1293 293 1309 327
rect 1377 293 1393 327
rect 1451 293 1467 327
rect 1535 293 1551 327
rect -1597 243 -1563 259
rect -1597 51 -1563 67
rect -1439 243 -1405 259
rect -1439 51 -1405 67
rect -1281 243 -1247 259
rect -1281 51 -1247 67
rect -1123 243 -1089 259
rect -1123 51 -1089 67
rect -965 243 -931 259
rect -965 51 -931 67
rect -807 243 -773 259
rect -807 51 -773 67
rect -649 243 -615 259
rect -649 51 -615 67
rect -491 243 -457 259
rect -491 51 -457 67
rect -333 243 -299 259
rect -333 51 -299 67
rect -175 243 -141 259
rect -175 51 -141 67
rect -17 243 17 259
rect -17 51 17 67
rect 141 243 175 259
rect 141 51 175 67
rect 299 243 333 259
rect 299 51 333 67
rect 457 243 491 259
rect 457 51 491 67
rect 615 243 649 259
rect 615 51 649 67
rect 773 243 807 259
rect 773 51 807 67
rect 931 243 965 259
rect 931 51 965 67
rect 1089 243 1123 259
rect 1089 51 1123 67
rect 1247 243 1281 259
rect 1247 51 1281 67
rect 1405 243 1439 259
rect 1405 51 1439 67
rect 1563 243 1597 259
rect 1563 51 1597 67
rect -1551 -17 -1535 17
rect -1467 -17 -1451 17
rect -1393 -17 -1377 17
rect -1309 -17 -1293 17
rect -1235 -17 -1219 17
rect -1151 -17 -1135 17
rect -1077 -17 -1061 17
rect -993 -17 -977 17
rect -919 -17 -903 17
rect -835 -17 -819 17
rect -761 -17 -745 17
rect -677 -17 -661 17
rect -603 -17 -587 17
rect -519 -17 -503 17
rect -445 -17 -429 17
rect -361 -17 -345 17
rect -287 -17 -271 17
rect -203 -17 -187 17
rect -129 -17 -113 17
rect -45 -17 -29 17
rect 29 -17 45 17
rect 113 -17 129 17
rect 187 -17 203 17
rect 271 -17 287 17
rect 345 -17 361 17
rect 429 -17 445 17
rect 503 -17 519 17
rect 587 -17 603 17
rect 661 -17 677 17
rect 745 -17 761 17
rect 819 -17 835 17
rect 903 -17 919 17
rect 977 -17 993 17
rect 1061 -17 1077 17
rect 1135 -17 1151 17
rect 1219 -17 1235 17
rect 1293 -17 1309 17
rect 1377 -17 1393 17
rect 1451 -17 1467 17
rect 1535 -17 1551 17
rect -1597 -67 -1563 -51
rect -1597 -259 -1563 -243
rect -1439 -67 -1405 -51
rect -1439 -259 -1405 -243
rect -1281 -67 -1247 -51
rect -1281 -259 -1247 -243
rect -1123 -67 -1089 -51
rect -1123 -259 -1089 -243
rect -965 -67 -931 -51
rect -965 -259 -931 -243
rect -807 -67 -773 -51
rect -807 -259 -773 -243
rect -649 -67 -615 -51
rect -649 -259 -615 -243
rect -491 -67 -457 -51
rect -491 -259 -457 -243
rect -333 -67 -299 -51
rect -333 -259 -299 -243
rect -175 -67 -141 -51
rect -175 -259 -141 -243
rect -17 -67 17 -51
rect -17 -259 17 -243
rect 141 -67 175 -51
rect 141 -259 175 -243
rect 299 -67 333 -51
rect 299 -259 333 -243
rect 457 -67 491 -51
rect 457 -259 491 -243
rect 615 -67 649 -51
rect 615 -259 649 -243
rect 773 -67 807 -51
rect 773 -259 807 -243
rect 931 -67 965 -51
rect 931 -259 965 -243
rect 1089 -67 1123 -51
rect 1089 -259 1123 -243
rect 1247 -67 1281 -51
rect 1247 -259 1281 -243
rect 1405 -67 1439 -51
rect 1405 -259 1439 -243
rect 1563 -67 1597 -51
rect 1563 -259 1597 -243
rect -1551 -327 -1535 -293
rect -1467 -327 -1451 -293
rect -1393 -327 -1377 -293
rect -1309 -327 -1293 -293
rect -1235 -327 -1219 -293
rect -1151 -327 -1135 -293
rect -1077 -327 -1061 -293
rect -993 -327 -977 -293
rect -919 -327 -903 -293
rect -835 -327 -819 -293
rect -761 -327 -745 -293
rect -677 -327 -661 -293
rect -603 -327 -587 -293
rect -519 -327 -503 -293
rect -445 -327 -429 -293
rect -361 -327 -345 -293
rect -287 -327 -271 -293
rect -203 -327 -187 -293
rect -129 -327 -113 -293
rect -45 -327 -29 -293
rect 29 -327 45 -293
rect 113 -327 129 -293
rect 187 -327 203 -293
rect 271 -327 287 -293
rect 345 -327 361 -293
rect 429 -327 445 -293
rect 503 -327 519 -293
rect 587 -327 603 -293
rect 661 -327 677 -293
rect 745 -327 761 -293
rect 819 -327 835 -293
rect 903 -327 919 -293
rect 977 -327 993 -293
rect 1061 -327 1077 -293
rect 1135 -327 1151 -293
rect 1219 -327 1235 -293
rect 1293 -327 1309 -293
rect 1377 -327 1393 -293
rect 1451 -327 1467 -293
rect 1535 -327 1551 -293
rect -1597 -377 -1563 -361
rect -1597 -569 -1563 -553
rect -1439 -377 -1405 -361
rect -1439 -569 -1405 -553
rect -1281 -377 -1247 -361
rect -1281 -569 -1247 -553
rect -1123 -377 -1089 -361
rect -1123 -569 -1089 -553
rect -965 -377 -931 -361
rect -965 -569 -931 -553
rect -807 -377 -773 -361
rect -807 -569 -773 -553
rect -649 -377 -615 -361
rect -649 -569 -615 -553
rect -491 -377 -457 -361
rect -491 -569 -457 -553
rect -333 -377 -299 -361
rect -333 -569 -299 -553
rect -175 -377 -141 -361
rect -175 -569 -141 -553
rect -17 -377 17 -361
rect -17 -569 17 -553
rect 141 -377 175 -361
rect 141 -569 175 -553
rect 299 -377 333 -361
rect 299 -569 333 -553
rect 457 -377 491 -361
rect 457 -569 491 -553
rect 615 -377 649 -361
rect 615 -569 649 -553
rect 773 -377 807 -361
rect 773 -569 807 -553
rect 931 -377 965 -361
rect 931 -569 965 -553
rect 1089 -377 1123 -361
rect 1089 -569 1123 -553
rect 1247 -377 1281 -361
rect 1247 -569 1281 -553
rect 1405 -377 1439 -361
rect 1405 -569 1439 -553
rect 1563 -377 1597 -361
rect 1563 -569 1597 -553
rect -1551 -637 -1535 -603
rect -1467 -637 -1451 -603
rect -1393 -637 -1377 -603
rect -1309 -637 -1293 -603
rect -1235 -637 -1219 -603
rect -1151 -637 -1135 -603
rect -1077 -637 -1061 -603
rect -993 -637 -977 -603
rect -919 -637 -903 -603
rect -835 -637 -819 -603
rect -761 -637 -745 -603
rect -677 -637 -661 -603
rect -603 -637 -587 -603
rect -519 -637 -503 -603
rect -445 -637 -429 -603
rect -361 -637 -345 -603
rect -287 -637 -271 -603
rect -203 -637 -187 -603
rect -129 -637 -113 -603
rect -45 -637 -29 -603
rect 29 -637 45 -603
rect 113 -637 129 -603
rect 187 -637 203 -603
rect 271 -637 287 -603
rect 345 -637 361 -603
rect 429 -637 445 -603
rect 503 -637 519 -603
rect 587 -637 603 -603
rect 661 -637 677 -603
rect 745 -637 761 -603
rect 819 -637 835 -603
rect 903 -637 919 -603
rect 977 -637 993 -603
rect 1061 -637 1077 -603
rect 1135 -637 1151 -603
rect 1219 -637 1235 -603
rect 1293 -637 1309 -603
rect 1377 -637 1393 -603
rect 1451 -637 1467 -603
rect 1535 -637 1551 -603
rect -1597 -687 -1563 -671
rect -1597 -879 -1563 -863
rect -1439 -687 -1405 -671
rect -1439 -879 -1405 -863
rect -1281 -687 -1247 -671
rect -1281 -879 -1247 -863
rect -1123 -687 -1089 -671
rect -1123 -879 -1089 -863
rect -965 -687 -931 -671
rect -965 -879 -931 -863
rect -807 -687 -773 -671
rect -807 -879 -773 -863
rect -649 -687 -615 -671
rect -649 -879 -615 -863
rect -491 -687 -457 -671
rect -491 -879 -457 -863
rect -333 -687 -299 -671
rect -333 -879 -299 -863
rect -175 -687 -141 -671
rect -175 -879 -141 -863
rect -17 -687 17 -671
rect -17 -879 17 -863
rect 141 -687 175 -671
rect 141 -879 175 -863
rect 299 -687 333 -671
rect 299 -879 333 -863
rect 457 -687 491 -671
rect 457 -879 491 -863
rect 615 -687 649 -671
rect 615 -879 649 -863
rect 773 -687 807 -671
rect 773 -879 807 -863
rect 931 -687 965 -671
rect 931 -879 965 -863
rect 1089 -687 1123 -671
rect 1089 -879 1123 -863
rect 1247 -687 1281 -671
rect 1247 -879 1281 -863
rect 1405 -687 1439 -671
rect 1405 -879 1439 -863
rect 1563 -687 1597 -671
rect 1563 -879 1597 -863
rect -1551 -947 -1535 -913
rect -1467 -947 -1451 -913
rect -1393 -947 -1377 -913
rect -1309 -947 -1293 -913
rect -1235 -947 -1219 -913
rect -1151 -947 -1135 -913
rect -1077 -947 -1061 -913
rect -993 -947 -977 -913
rect -919 -947 -903 -913
rect -835 -947 -819 -913
rect -761 -947 -745 -913
rect -677 -947 -661 -913
rect -603 -947 -587 -913
rect -519 -947 -503 -913
rect -445 -947 -429 -913
rect -361 -947 -345 -913
rect -287 -947 -271 -913
rect -203 -947 -187 -913
rect -129 -947 -113 -913
rect -45 -947 -29 -913
rect 29 -947 45 -913
rect 113 -947 129 -913
rect 187 -947 203 -913
rect 271 -947 287 -913
rect 345 -947 361 -913
rect 429 -947 445 -913
rect 503 -947 519 -913
rect 587 -947 603 -913
rect 661 -947 677 -913
rect 745 -947 761 -913
rect 819 -947 835 -913
rect 903 -947 919 -913
rect 977 -947 993 -913
rect 1061 -947 1077 -913
rect 1135 -947 1151 -913
rect 1219 -947 1235 -913
rect 1293 -947 1309 -913
rect 1377 -947 1393 -913
rect 1451 -947 1467 -913
rect 1535 -947 1551 -913
rect -1597 -997 -1563 -981
rect -1597 -1189 -1563 -1173
rect -1439 -997 -1405 -981
rect -1439 -1189 -1405 -1173
rect -1281 -997 -1247 -981
rect -1281 -1189 -1247 -1173
rect -1123 -997 -1089 -981
rect -1123 -1189 -1089 -1173
rect -965 -997 -931 -981
rect -965 -1189 -931 -1173
rect -807 -997 -773 -981
rect -807 -1189 -773 -1173
rect -649 -997 -615 -981
rect -649 -1189 -615 -1173
rect -491 -997 -457 -981
rect -491 -1189 -457 -1173
rect -333 -997 -299 -981
rect -333 -1189 -299 -1173
rect -175 -997 -141 -981
rect -175 -1189 -141 -1173
rect -17 -997 17 -981
rect -17 -1189 17 -1173
rect 141 -997 175 -981
rect 141 -1189 175 -1173
rect 299 -997 333 -981
rect 299 -1189 333 -1173
rect 457 -997 491 -981
rect 457 -1189 491 -1173
rect 615 -997 649 -981
rect 615 -1189 649 -1173
rect 773 -997 807 -981
rect 773 -1189 807 -1173
rect 931 -997 965 -981
rect 931 -1189 965 -1173
rect 1089 -997 1123 -981
rect 1089 -1189 1123 -1173
rect 1247 -997 1281 -981
rect 1247 -1189 1281 -1173
rect 1405 -997 1439 -981
rect 1405 -1189 1439 -1173
rect 1563 -997 1597 -981
rect 1563 -1189 1597 -1173
rect -1551 -1257 -1535 -1223
rect -1467 -1257 -1451 -1223
rect -1393 -1257 -1377 -1223
rect -1309 -1257 -1293 -1223
rect -1235 -1257 -1219 -1223
rect -1151 -1257 -1135 -1223
rect -1077 -1257 -1061 -1223
rect -993 -1257 -977 -1223
rect -919 -1257 -903 -1223
rect -835 -1257 -819 -1223
rect -761 -1257 -745 -1223
rect -677 -1257 -661 -1223
rect -603 -1257 -587 -1223
rect -519 -1257 -503 -1223
rect -445 -1257 -429 -1223
rect -361 -1257 -345 -1223
rect -287 -1257 -271 -1223
rect -203 -1257 -187 -1223
rect -129 -1257 -113 -1223
rect -45 -1257 -29 -1223
rect 29 -1257 45 -1223
rect 113 -1257 129 -1223
rect 187 -1257 203 -1223
rect 271 -1257 287 -1223
rect 345 -1257 361 -1223
rect 429 -1257 445 -1223
rect 503 -1257 519 -1223
rect 587 -1257 603 -1223
rect 661 -1257 677 -1223
rect 745 -1257 761 -1223
rect 819 -1257 835 -1223
rect 903 -1257 919 -1223
rect 977 -1257 993 -1223
rect 1061 -1257 1077 -1223
rect 1135 -1257 1151 -1223
rect 1219 -1257 1235 -1223
rect 1293 -1257 1309 -1223
rect 1377 -1257 1393 -1223
rect 1451 -1257 1467 -1223
rect 1535 -1257 1551 -1223
rect -1597 -1307 -1563 -1291
rect -1597 -1499 -1563 -1483
rect -1439 -1307 -1405 -1291
rect -1439 -1499 -1405 -1483
rect -1281 -1307 -1247 -1291
rect -1281 -1499 -1247 -1483
rect -1123 -1307 -1089 -1291
rect -1123 -1499 -1089 -1483
rect -965 -1307 -931 -1291
rect -965 -1499 -931 -1483
rect -807 -1307 -773 -1291
rect -807 -1499 -773 -1483
rect -649 -1307 -615 -1291
rect -649 -1499 -615 -1483
rect -491 -1307 -457 -1291
rect -491 -1499 -457 -1483
rect -333 -1307 -299 -1291
rect -333 -1499 -299 -1483
rect -175 -1307 -141 -1291
rect -175 -1499 -141 -1483
rect -17 -1307 17 -1291
rect -17 -1499 17 -1483
rect 141 -1307 175 -1291
rect 141 -1499 175 -1483
rect 299 -1307 333 -1291
rect 299 -1499 333 -1483
rect 457 -1307 491 -1291
rect 457 -1499 491 -1483
rect 615 -1307 649 -1291
rect 615 -1499 649 -1483
rect 773 -1307 807 -1291
rect 773 -1499 807 -1483
rect 931 -1307 965 -1291
rect 931 -1499 965 -1483
rect 1089 -1307 1123 -1291
rect 1089 -1499 1123 -1483
rect 1247 -1307 1281 -1291
rect 1247 -1499 1281 -1483
rect 1405 -1307 1439 -1291
rect 1405 -1499 1439 -1483
rect 1563 -1307 1597 -1291
rect 1563 -1499 1597 -1483
rect -1551 -1567 -1535 -1533
rect -1467 -1567 -1451 -1533
rect -1393 -1567 -1377 -1533
rect -1309 -1567 -1293 -1533
rect -1235 -1567 -1219 -1533
rect -1151 -1567 -1135 -1533
rect -1077 -1567 -1061 -1533
rect -993 -1567 -977 -1533
rect -919 -1567 -903 -1533
rect -835 -1567 -819 -1533
rect -761 -1567 -745 -1533
rect -677 -1567 -661 -1533
rect -603 -1567 -587 -1533
rect -519 -1567 -503 -1533
rect -445 -1567 -429 -1533
rect -361 -1567 -345 -1533
rect -287 -1567 -271 -1533
rect -203 -1567 -187 -1533
rect -129 -1567 -113 -1533
rect -45 -1567 -29 -1533
rect 29 -1567 45 -1533
rect 113 -1567 129 -1533
rect 187 -1567 203 -1533
rect 271 -1567 287 -1533
rect 345 -1567 361 -1533
rect 429 -1567 445 -1533
rect 503 -1567 519 -1533
rect 587 -1567 603 -1533
rect 661 -1567 677 -1533
rect 745 -1567 761 -1533
rect 819 -1567 835 -1533
rect 903 -1567 919 -1533
rect 977 -1567 993 -1533
rect 1061 -1567 1077 -1533
rect 1135 -1567 1151 -1533
rect 1219 -1567 1235 -1533
rect 1293 -1567 1309 -1533
rect 1377 -1567 1393 -1533
rect 1451 -1567 1467 -1533
rect 1535 -1567 1551 -1533
rect -1731 -1671 -1697 -1609
rect 1697 -1671 1731 -1609
rect -1731 -1705 -1635 -1671
rect 1635 -1705 1731 -1671
<< viali >>
rect -1535 1533 -1467 1567
rect -1377 1533 -1309 1567
rect -1219 1533 -1151 1567
rect -1061 1533 -993 1567
rect -903 1533 -835 1567
rect -745 1533 -677 1567
rect -587 1533 -519 1567
rect -429 1533 -361 1567
rect -271 1533 -203 1567
rect -113 1533 -45 1567
rect 45 1533 113 1567
rect 203 1533 271 1567
rect 361 1533 429 1567
rect 519 1533 587 1567
rect 677 1533 745 1567
rect 835 1533 903 1567
rect 993 1533 1061 1567
rect 1151 1533 1219 1567
rect 1309 1533 1377 1567
rect 1467 1533 1535 1567
rect -1597 1307 -1563 1483
rect -1439 1307 -1405 1483
rect -1281 1307 -1247 1483
rect -1123 1307 -1089 1483
rect -965 1307 -931 1483
rect -807 1307 -773 1483
rect -649 1307 -615 1483
rect -491 1307 -457 1483
rect -333 1307 -299 1483
rect -175 1307 -141 1483
rect -17 1307 17 1483
rect 141 1307 175 1483
rect 299 1307 333 1483
rect 457 1307 491 1483
rect 615 1307 649 1483
rect 773 1307 807 1483
rect 931 1307 965 1483
rect 1089 1307 1123 1483
rect 1247 1307 1281 1483
rect 1405 1307 1439 1483
rect 1563 1307 1597 1483
rect -1535 1223 -1467 1257
rect -1377 1223 -1309 1257
rect -1219 1223 -1151 1257
rect -1061 1223 -993 1257
rect -903 1223 -835 1257
rect -745 1223 -677 1257
rect -587 1223 -519 1257
rect -429 1223 -361 1257
rect -271 1223 -203 1257
rect -113 1223 -45 1257
rect 45 1223 113 1257
rect 203 1223 271 1257
rect 361 1223 429 1257
rect 519 1223 587 1257
rect 677 1223 745 1257
rect 835 1223 903 1257
rect 993 1223 1061 1257
rect 1151 1223 1219 1257
rect 1309 1223 1377 1257
rect 1467 1223 1535 1257
rect -1597 997 -1563 1173
rect -1439 997 -1405 1173
rect -1281 997 -1247 1173
rect -1123 997 -1089 1173
rect -965 997 -931 1173
rect -807 997 -773 1173
rect -649 997 -615 1173
rect -491 997 -457 1173
rect -333 997 -299 1173
rect -175 997 -141 1173
rect -17 997 17 1173
rect 141 997 175 1173
rect 299 997 333 1173
rect 457 997 491 1173
rect 615 997 649 1173
rect 773 997 807 1173
rect 931 997 965 1173
rect 1089 997 1123 1173
rect 1247 997 1281 1173
rect 1405 997 1439 1173
rect 1563 997 1597 1173
rect -1535 913 -1467 947
rect -1377 913 -1309 947
rect -1219 913 -1151 947
rect -1061 913 -993 947
rect -903 913 -835 947
rect -745 913 -677 947
rect -587 913 -519 947
rect -429 913 -361 947
rect -271 913 -203 947
rect -113 913 -45 947
rect 45 913 113 947
rect 203 913 271 947
rect 361 913 429 947
rect 519 913 587 947
rect 677 913 745 947
rect 835 913 903 947
rect 993 913 1061 947
rect 1151 913 1219 947
rect 1309 913 1377 947
rect 1467 913 1535 947
rect -1597 687 -1563 863
rect -1439 687 -1405 863
rect -1281 687 -1247 863
rect -1123 687 -1089 863
rect -965 687 -931 863
rect -807 687 -773 863
rect -649 687 -615 863
rect -491 687 -457 863
rect -333 687 -299 863
rect -175 687 -141 863
rect -17 687 17 863
rect 141 687 175 863
rect 299 687 333 863
rect 457 687 491 863
rect 615 687 649 863
rect 773 687 807 863
rect 931 687 965 863
rect 1089 687 1123 863
rect 1247 687 1281 863
rect 1405 687 1439 863
rect 1563 687 1597 863
rect -1535 603 -1467 637
rect -1377 603 -1309 637
rect -1219 603 -1151 637
rect -1061 603 -993 637
rect -903 603 -835 637
rect -745 603 -677 637
rect -587 603 -519 637
rect -429 603 -361 637
rect -271 603 -203 637
rect -113 603 -45 637
rect 45 603 113 637
rect 203 603 271 637
rect 361 603 429 637
rect 519 603 587 637
rect 677 603 745 637
rect 835 603 903 637
rect 993 603 1061 637
rect 1151 603 1219 637
rect 1309 603 1377 637
rect 1467 603 1535 637
rect -1597 377 -1563 553
rect -1439 377 -1405 553
rect -1281 377 -1247 553
rect -1123 377 -1089 553
rect -965 377 -931 553
rect -807 377 -773 553
rect -649 377 -615 553
rect -491 377 -457 553
rect -333 377 -299 553
rect -175 377 -141 553
rect -17 377 17 553
rect 141 377 175 553
rect 299 377 333 553
rect 457 377 491 553
rect 615 377 649 553
rect 773 377 807 553
rect 931 377 965 553
rect 1089 377 1123 553
rect 1247 377 1281 553
rect 1405 377 1439 553
rect 1563 377 1597 553
rect -1535 293 -1467 327
rect -1377 293 -1309 327
rect -1219 293 -1151 327
rect -1061 293 -993 327
rect -903 293 -835 327
rect -745 293 -677 327
rect -587 293 -519 327
rect -429 293 -361 327
rect -271 293 -203 327
rect -113 293 -45 327
rect 45 293 113 327
rect 203 293 271 327
rect 361 293 429 327
rect 519 293 587 327
rect 677 293 745 327
rect 835 293 903 327
rect 993 293 1061 327
rect 1151 293 1219 327
rect 1309 293 1377 327
rect 1467 293 1535 327
rect -1597 67 -1563 243
rect -1439 67 -1405 243
rect -1281 67 -1247 243
rect -1123 67 -1089 243
rect -965 67 -931 243
rect -807 67 -773 243
rect -649 67 -615 243
rect -491 67 -457 243
rect -333 67 -299 243
rect -175 67 -141 243
rect -17 67 17 243
rect 141 67 175 243
rect 299 67 333 243
rect 457 67 491 243
rect 615 67 649 243
rect 773 67 807 243
rect 931 67 965 243
rect 1089 67 1123 243
rect 1247 67 1281 243
rect 1405 67 1439 243
rect 1563 67 1597 243
rect -1535 -17 -1467 17
rect -1377 -17 -1309 17
rect -1219 -17 -1151 17
rect -1061 -17 -993 17
rect -903 -17 -835 17
rect -745 -17 -677 17
rect -587 -17 -519 17
rect -429 -17 -361 17
rect -271 -17 -203 17
rect -113 -17 -45 17
rect 45 -17 113 17
rect 203 -17 271 17
rect 361 -17 429 17
rect 519 -17 587 17
rect 677 -17 745 17
rect 835 -17 903 17
rect 993 -17 1061 17
rect 1151 -17 1219 17
rect 1309 -17 1377 17
rect 1467 -17 1535 17
rect -1597 -243 -1563 -67
rect -1439 -243 -1405 -67
rect -1281 -243 -1247 -67
rect -1123 -243 -1089 -67
rect -965 -243 -931 -67
rect -807 -243 -773 -67
rect -649 -243 -615 -67
rect -491 -243 -457 -67
rect -333 -243 -299 -67
rect -175 -243 -141 -67
rect -17 -243 17 -67
rect 141 -243 175 -67
rect 299 -243 333 -67
rect 457 -243 491 -67
rect 615 -243 649 -67
rect 773 -243 807 -67
rect 931 -243 965 -67
rect 1089 -243 1123 -67
rect 1247 -243 1281 -67
rect 1405 -243 1439 -67
rect 1563 -243 1597 -67
rect -1535 -327 -1467 -293
rect -1377 -327 -1309 -293
rect -1219 -327 -1151 -293
rect -1061 -327 -993 -293
rect -903 -327 -835 -293
rect -745 -327 -677 -293
rect -587 -327 -519 -293
rect -429 -327 -361 -293
rect -271 -327 -203 -293
rect -113 -327 -45 -293
rect 45 -327 113 -293
rect 203 -327 271 -293
rect 361 -327 429 -293
rect 519 -327 587 -293
rect 677 -327 745 -293
rect 835 -327 903 -293
rect 993 -327 1061 -293
rect 1151 -327 1219 -293
rect 1309 -327 1377 -293
rect 1467 -327 1535 -293
rect -1597 -553 -1563 -377
rect -1439 -553 -1405 -377
rect -1281 -553 -1247 -377
rect -1123 -553 -1089 -377
rect -965 -553 -931 -377
rect -807 -553 -773 -377
rect -649 -553 -615 -377
rect -491 -553 -457 -377
rect -333 -553 -299 -377
rect -175 -553 -141 -377
rect -17 -553 17 -377
rect 141 -553 175 -377
rect 299 -553 333 -377
rect 457 -553 491 -377
rect 615 -553 649 -377
rect 773 -553 807 -377
rect 931 -553 965 -377
rect 1089 -553 1123 -377
rect 1247 -553 1281 -377
rect 1405 -553 1439 -377
rect 1563 -553 1597 -377
rect -1535 -637 -1467 -603
rect -1377 -637 -1309 -603
rect -1219 -637 -1151 -603
rect -1061 -637 -993 -603
rect -903 -637 -835 -603
rect -745 -637 -677 -603
rect -587 -637 -519 -603
rect -429 -637 -361 -603
rect -271 -637 -203 -603
rect -113 -637 -45 -603
rect 45 -637 113 -603
rect 203 -637 271 -603
rect 361 -637 429 -603
rect 519 -637 587 -603
rect 677 -637 745 -603
rect 835 -637 903 -603
rect 993 -637 1061 -603
rect 1151 -637 1219 -603
rect 1309 -637 1377 -603
rect 1467 -637 1535 -603
rect -1597 -863 -1563 -687
rect -1439 -863 -1405 -687
rect -1281 -863 -1247 -687
rect -1123 -863 -1089 -687
rect -965 -863 -931 -687
rect -807 -863 -773 -687
rect -649 -863 -615 -687
rect -491 -863 -457 -687
rect -333 -863 -299 -687
rect -175 -863 -141 -687
rect -17 -863 17 -687
rect 141 -863 175 -687
rect 299 -863 333 -687
rect 457 -863 491 -687
rect 615 -863 649 -687
rect 773 -863 807 -687
rect 931 -863 965 -687
rect 1089 -863 1123 -687
rect 1247 -863 1281 -687
rect 1405 -863 1439 -687
rect 1563 -863 1597 -687
rect -1535 -947 -1467 -913
rect -1377 -947 -1309 -913
rect -1219 -947 -1151 -913
rect -1061 -947 -993 -913
rect -903 -947 -835 -913
rect -745 -947 -677 -913
rect -587 -947 -519 -913
rect -429 -947 -361 -913
rect -271 -947 -203 -913
rect -113 -947 -45 -913
rect 45 -947 113 -913
rect 203 -947 271 -913
rect 361 -947 429 -913
rect 519 -947 587 -913
rect 677 -947 745 -913
rect 835 -947 903 -913
rect 993 -947 1061 -913
rect 1151 -947 1219 -913
rect 1309 -947 1377 -913
rect 1467 -947 1535 -913
rect -1597 -1173 -1563 -997
rect -1439 -1173 -1405 -997
rect -1281 -1173 -1247 -997
rect -1123 -1173 -1089 -997
rect -965 -1173 -931 -997
rect -807 -1173 -773 -997
rect -649 -1173 -615 -997
rect -491 -1173 -457 -997
rect -333 -1173 -299 -997
rect -175 -1173 -141 -997
rect -17 -1173 17 -997
rect 141 -1173 175 -997
rect 299 -1173 333 -997
rect 457 -1173 491 -997
rect 615 -1173 649 -997
rect 773 -1173 807 -997
rect 931 -1173 965 -997
rect 1089 -1173 1123 -997
rect 1247 -1173 1281 -997
rect 1405 -1173 1439 -997
rect 1563 -1173 1597 -997
rect -1535 -1257 -1467 -1223
rect -1377 -1257 -1309 -1223
rect -1219 -1257 -1151 -1223
rect -1061 -1257 -993 -1223
rect -903 -1257 -835 -1223
rect -745 -1257 -677 -1223
rect -587 -1257 -519 -1223
rect -429 -1257 -361 -1223
rect -271 -1257 -203 -1223
rect -113 -1257 -45 -1223
rect 45 -1257 113 -1223
rect 203 -1257 271 -1223
rect 361 -1257 429 -1223
rect 519 -1257 587 -1223
rect 677 -1257 745 -1223
rect 835 -1257 903 -1223
rect 993 -1257 1061 -1223
rect 1151 -1257 1219 -1223
rect 1309 -1257 1377 -1223
rect 1467 -1257 1535 -1223
rect -1597 -1483 -1563 -1307
rect -1439 -1483 -1405 -1307
rect -1281 -1483 -1247 -1307
rect -1123 -1483 -1089 -1307
rect -965 -1483 -931 -1307
rect -807 -1483 -773 -1307
rect -649 -1483 -615 -1307
rect -491 -1483 -457 -1307
rect -333 -1483 -299 -1307
rect -175 -1483 -141 -1307
rect -17 -1483 17 -1307
rect 141 -1483 175 -1307
rect 299 -1483 333 -1307
rect 457 -1483 491 -1307
rect 615 -1483 649 -1307
rect 773 -1483 807 -1307
rect 931 -1483 965 -1307
rect 1089 -1483 1123 -1307
rect 1247 -1483 1281 -1307
rect 1405 -1483 1439 -1307
rect 1563 -1483 1597 -1307
rect -1535 -1567 -1467 -1533
rect -1377 -1567 -1309 -1533
rect -1219 -1567 -1151 -1533
rect -1061 -1567 -993 -1533
rect -903 -1567 -835 -1533
rect -745 -1567 -677 -1533
rect -587 -1567 -519 -1533
rect -429 -1567 -361 -1533
rect -271 -1567 -203 -1533
rect -113 -1567 -45 -1533
rect 45 -1567 113 -1533
rect 203 -1567 271 -1533
rect 361 -1567 429 -1533
rect 519 -1567 587 -1533
rect 677 -1567 745 -1533
rect 835 -1567 903 -1533
rect 993 -1567 1061 -1533
rect 1151 -1567 1219 -1533
rect 1309 -1567 1377 -1533
rect 1467 -1567 1535 -1533
<< metal1 >>
rect -1547 1567 -1455 1573
rect -1547 1533 -1535 1567
rect -1467 1533 -1455 1567
rect -1547 1527 -1455 1533
rect -1389 1567 -1297 1573
rect -1389 1533 -1377 1567
rect -1309 1533 -1297 1567
rect -1389 1527 -1297 1533
rect -1231 1567 -1139 1573
rect -1231 1533 -1219 1567
rect -1151 1533 -1139 1567
rect -1231 1527 -1139 1533
rect -1073 1567 -981 1573
rect -1073 1533 -1061 1567
rect -993 1533 -981 1567
rect -1073 1527 -981 1533
rect -915 1567 -823 1573
rect -915 1533 -903 1567
rect -835 1533 -823 1567
rect -915 1527 -823 1533
rect -757 1567 -665 1573
rect -757 1533 -745 1567
rect -677 1533 -665 1567
rect -757 1527 -665 1533
rect -599 1567 -507 1573
rect -599 1533 -587 1567
rect -519 1533 -507 1567
rect -599 1527 -507 1533
rect -441 1567 -349 1573
rect -441 1533 -429 1567
rect -361 1533 -349 1567
rect -441 1527 -349 1533
rect -283 1567 -191 1573
rect -283 1533 -271 1567
rect -203 1533 -191 1567
rect -283 1527 -191 1533
rect -125 1567 -33 1573
rect -125 1533 -113 1567
rect -45 1533 -33 1567
rect -125 1527 -33 1533
rect 33 1567 125 1573
rect 33 1533 45 1567
rect 113 1533 125 1567
rect 33 1527 125 1533
rect 191 1567 283 1573
rect 191 1533 203 1567
rect 271 1533 283 1567
rect 191 1527 283 1533
rect 349 1567 441 1573
rect 349 1533 361 1567
rect 429 1533 441 1567
rect 349 1527 441 1533
rect 507 1567 599 1573
rect 507 1533 519 1567
rect 587 1533 599 1567
rect 507 1527 599 1533
rect 665 1567 757 1573
rect 665 1533 677 1567
rect 745 1533 757 1567
rect 665 1527 757 1533
rect 823 1567 915 1573
rect 823 1533 835 1567
rect 903 1533 915 1567
rect 823 1527 915 1533
rect 981 1567 1073 1573
rect 981 1533 993 1567
rect 1061 1533 1073 1567
rect 981 1527 1073 1533
rect 1139 1567 1231 1573
rect 1139 1533 1151 1567
rect 1219 1533 1231 1567
rect 1139 1527 1231 1533
rect 1297 1567 1389 1573
rect 1297 1533 1309 1567
rect 1377 1533 1389 1567
rect 1297 1527 1389 1533
rect 1455 1567 1547 1573
rect 1455 1533 1467 1567
rect 1535 1533 1547 1567
rect 1455 1527 1547 1533
rect -1603 1483 -1557 1495
rect -1603 1307 -1597 1483
rect -1563 1307 -1557 1483
rect -1603 1295 -1557 1307
rect -1445 1483 -1399 1495
rect -1445 1307 -1439 1483
rect -1405 1307 -1399 1483
rect -1445 1295 -1399 1307
rect -1287 1483 -1241 1495
rect -1287 1307 -1281 1483
rect -1247 1307 -1241 1483
rect -1287 1295 -1241 1307
rect -1129 1483 -1083 1495
rect -1129 1307 -1123 1483
rect -1089 1307 -1083 1483
rect -1129 1295 -1083 1307
rect -971 1483 -925 1495
rect -971 1307 -965 1483
rect -931 1307 -925 1483
rect -971 1295 -925 1307
rect -813 1483 -767 1495
rect -813 1307 -807 1483
rect -773 1307 -767 1483
rect -813 1295 -767 1307
rect -655 1483 -609 1495
rect -655 1307 -649 1483
rect -615 1307 -609 1483
rect -655 1295 -609 1307
rect -497 1483 -451 1495
rect -497 1307 -491 1483
rect -457 1307 -451 1483
rect -497 1295 -451 1307
rect -339 1483 -293 1495
rect -339 1307 -333 1483
rect -299 1307 -293 1483
rect -339 1295 -293 1307
rect -181 1483 -135 1495
rect -181 1307 -175 1483
rect -141 1307 -135 1483
rect -181 1295 -135 1307
rect -23 1483 23 1495
rect -23 1307 -17 1483
rect 17 1307 23 1483
rect -23 1295 23 1307
rect 135 1483 181 1495
rect 135 1307 141 1483
rect 175 1307 181 1483
rect 135 1295 181 1307
rect 293 1483 339 1495
rect 293 1307 299 1483
rect 333 1307 339 1483
rect 293 1295 339 1307
rect 451 1483 497 1495
rect 451 1307 457 1483
rect 491 1307 497 1483
rect 451 1295 497 1307
rect 609 1483 655 1495
rect 609 1307 615 1483
rect 649 1307 655 1483
rect 609 1295 655 1307
rect 767 1483 813 1495
rect 767 1307 773 1483
rect 807 1307 813 1483
rect 767 1295 813 1307
rect 925 1483 971 1495
rect 925 1307 931 1483
rect 965 1307 971 1483
rect 925 1295 971 1307
rect 1083 1483 1129 1495
rect 1083 1307 1089 1483
rect 1123 1307 1129 1483
rect 1083 1295 1129 1307
rect 1241 1483 1287 1495
rect 1241 1307 1247 1483
rect 1281 1307 1287 1483
rect 1241 1295 1287 1307
rect 1399 1483 1445 1495
rect 1399 1307 1405 1483
rect 1439 1307 1445 1483
rect 1399 1295 1445 1307
rect 1557 1483 1603 1495
rect 1557 1307 1563 1483
rect 1597 1307 1603 1483
rect 1557 1295 1603 1307
rect -1547 1257 -1455 1263
rect -1547 1223 -1535 1257
rect -1467 1223 -1455 1257
rect -1547 1217 -1455 1223
rect -1389 1257 -1297 1263
rect -1389 1223 -1377 1257
rect -1309 1223 -1297 1257
rect -1389 1217 -1297 1223
rect -1231 1257 -1139 1263
rect -1231 1223 -1219 1257
rect -1151 1223 -1139 1257
rect -1231 1217 -1139 1223
rect -1073 1257 -981 1263
rect -1073 1223 -1061 1257
rect -993 1223 -981 1257
rect -1073 1217 -981 1223
rect -915 1257 -823 1263
rect -915 1223 -903 1257
rect -835 1223 -823 1257
rect -915 1217 -823 1223
rect -757 1257 -665 1263
rect -757 1223 -745 1257
rect -677 1223 -665 1257
rect -757 1217 -665 1223
rect -599 1257 -507 1263
rect -599 1223 -587 1257
rect -519 1223 -507 1257
rect -599 1217 -507 1223
rect -441 1257 -349 1263
rect -441 1223 -429 1257
rect -361 1223 -349 1257
rect -441 1217 -349 1223
rect -283 1257 -191 1263
rect -283 1223 -271 1257
rect -203 1223 -191 1257
rect -283 1217 -191 1223
rect -125 1257 -33 1263
rect -125 1223 -113 1257
rect -45 1223 -33 1257
rect -125 1217 -33 1223
rect 33 1257 125 1263
rect 33 1223 45 1257
rect 113 1223 125 1257
rect 33 1217 125 1223
rect 191 1257 283 1263
rect 191 1223 203 1257
rect 271 1223 283 1257
rect 191 1217 283 1223
rect 349 1257 441 1263
rect 349 1223 361 1257
rect 429 1223 441 1257
rect 349 1217 441 1223
rect 507 1257 599 1263
rect 507 1223 519 1257
rect 587 1223 599 1257
rect 507 1217 599 1223
rect 665 1257 757 1263
rect 665 1223 677 1257
rect 745 1223 757 1257
rect 665 1217 757 1223
rect 823 1257 915 1263
rect 823 1223 835 1257
rect 903 1223 915 1257
rect 823 1217 915 1223
rect 981 1257 1073 1263
rect 981 1223 993 1257
rect 1061 1223 1073 1257
rect 981 1217 1073 1223
rect 1139 1257 1231 1263
rect 1139 1223 1151 1257
rect 1219 1223 1231 1257
rect 1139 1217 1231 1223
rect 1297 1257 1389 1263
rect 1297 1223 1309 1257
rect 1377 1223 1389 1257
rect 1297 1217 1389 1223
rect 1455 1257 1547 1263
rect 1455 1223 1467 1257
rect 1535 1223 1547 1257
rect 1455 1217 1547 1223
rect -1603 1173 -1557 1185
rect -1603 997 -1597 1173
rect -1563 997 -1557 1173
rect -1603 985 -1557 997
rect -1445 1173 -1399 1185
rect -1445 997 -1439 1173
rect -1405 997 -1399 1173
rect -1445 985 -1399 997
rect -1287 1173 -1241 1185
rect -1287 997 -1281 1173
rect -1247 997 -1241 1173
rect -1287 985 -1241 997
rect -1129 1173 -1083 1185
rect -1129 997 -1123 1173
rect -1089 997 -1083 1173
rect -1129 985 -1083 997
rect -971 1173 -925 1185
rect -971 997 -965 1173
rect -931 997 -925 1173
rect -971 985 -925 997
rect -813 1173 -767 1185
rect -813 997 -807 1173
rect -773 997 -767 1173
rect -813 985 -767 997
rect -655 1173 -609 1185
rect -655 997 -649 1173
rect -615 997 -609 1173
rect -655 985 -609 997
rect -497 1173 -451 1185
rect -497 997 -491 1173
rect -457 997 -451 1173
rect -497 985 -451 997
rect -339 1173 -293 1185
rect -339 997 -333 1173
rect -299 997 -293 1173
rect -339 985 -293 997
rect -181 1173 -135 1185
rect -181 997 -175 1173
rect -141 997 -135 1173
rect -181 985 -135 997
rect -23 1173 23 1185
rect -23 997 -17 1173
rect 17 997 23 1173
rect -23 985 23 997
rect 135 1173 181 1185
rect 135 997 141 1173
rect 175 997 181 1173
rect 135 985 181 997
rect 293 1173 339 1185
rect 293 997 299 1173
rect 333 997 339 1173
rect 293 985 339 997
rect 451 1173 497 1185
rect 451 997 457 1173
rect 491 997 497 1173
rect 451 985 497 997
rect 609 1173 655 1185
rect 609 997 615 1173
rect 649 997 655 1173
rect 609 985 655 997
rect 767 1173 813 1185
rect 767 997 773 1173
rect 807 997 813 1173
rect 767 985 813 997
rect 925 1173 971 1185
rect 925 997 931 1173
rect 965 997 971 1173
rect 925 985 971 997
rect 1083 1173 1129 1185
rect 1083 997 1089 1173
rect 1123 997 1129 1173
rect 1083 985 1129 997
rect 1241 1173 1287 1185
rect 1241 997 1247 1173
rect 1281 997 1287 1173
rect 1241 985 1287 997
rect 1399 1173 1445 1185
rect 1399 997 1405 1173
rect 1439 997 1445 1173
rect 1399 985 1445 997
rect 1557 1173 1603 1185
rect 1557 997 1563 1173
rect 1597 997 1603 1173
rect 1557 985 1603 997
rect -1547 947 -1455 953
rect -1547 913 -1535 947
rect -1467 913 -1455 947
rect -1547 907 -1455 913
rect -1389 947 -1297 953
rect -1389 913 -1377 947
rect -1309 913 -1297 947
rect -1389 907 -1297 913
rect -1231 947 -1139 953
rect -1231 913 -1219 947
rect -1151 913 -1139 947
rect -1231 907 -1139 913
rect -1073 947 -981 953
rect -1073 913 -1061 947
rect -993 913 -981 947
rect -1073 907 -981 913
rect -915 947 -823 953
rect -915 913 -903 947
rect -835 913 -823 947
rect -915 907 -823 913
rect -757 947 -665 953
rect -757 913 -745 947
rect -677 913 -665 947
rect -757 907 -665 913
rect -599 947 -507 953
rect -599 913 -587 947
rect -519 913 -507 947
rect -599 907 -507 913
rect -441 947 -349 953
rect -441 913 -429 947
rect -361 913 -349 947
rect -441 907 -349 913
rect -283 947 -191 953
rect -283 913 -271 947
rect -203 913 -191 947
rect -283 907 -191 913
rect -125 947 -33 953
rect -125 913 -113 947
rect -45 913 -33 947
rect -125 907 -33 913
rect 33 947 125 953
rect 33 913 45 947
rect 113 913 125 947
rect 33 907 125 913
rect 191 947 283 953
rect 191 913 203 947
rect 271 913 283 947
rect 191 907 283 913
rect 349 947 441 953
rect 349 913 361 947
rect 429 913 441 947
rect 349 907 441 913
rect 507 947 599 953
rect 507 913 519 947
rect 587 913 599 947
rect 507 907 599 913
rect 665 947 757 953
rect 665 913 677 947
rect 745 913 757 947
rect 665 907 757 913
rect 823 947 915 953
rect 823 913 835 947
rect 903 913 915 947
rect 823 907 915 913
rect 981 947 1073 953
rect 981 913 993 947
rect 1061 913 1073 947
rect 981 907 1073 913
rect 1139 947 1231 953
rect 1139 913 1151 947
rect 1219 913 1231 947
rect 1139 907 1231 913
rect 1297 947 1389 953
rect 1297 913 1309 947
rect 1377 913 1389 947
rect 1297 907 1389 913
rect 1455 947 1547 953
rect 1455 913 1467 947
rect 1535 913 1547 947
rect 1455 907 1547 913
rect -1603 863 -1557 875
rect -1603 687 -1597 863
rect -1563 687 -1557 863
rect -1603 675 -1557 687
rect -1445 863 -1399 875
rect -1445 687 -1439 863
rect -1405 687 -1399 863
rect -1445 675 -1399 687
rect -1287 863 -1241 875
rect -1287 687 -1281 863
rect -1247 687 -1241 863
rect -1287 675 -1241 687
rect -1129 863 -1083 875
rect -1129 687 -1123 863
rect -1089 687 -1083 863
rect -1129 675 -1083 687
rect -971 863 -925 875
rect -971 687 -965 863
rect -931 687 -925 863
rect -971 675 -925 687
rect -813 863 -767 875
rect -813 687 -807 863
rect -773 687 -767 863
rect -813 675 -767 687
rect -655 863 -609 875
rect -655 687 -649 863
rect -615 687 -609 863
rect -655 675 -609 687
rect -497 863 -451 875
rect -497 687 -491 863
rect -457 687 -451 863
rect -497 675 -451 687
rect -339 863 -293 875
rect -339 687 -333 863
rect -299 687 -293 863
rect -339 675 -293 687
rect -181 863 -135 875
rect -181 687 -175 863
rect -141 687 -135 863
rect -181 675 -135 687
rect -23 863 23 875
rect -23 687 -17 863
rect 17 687 23 863
rect -23 675 23 687
rect 135 863 181 875
rect 135 687 141 863
rect 175 687 181 863
rect 135 675 181 687
rect 293 863 339 875
rect 293 687 299 863
rect 333 687 339 863
rect 293 675 339 687
rect 451 863 497 875
rect 451 687 457 863
rect 491 687 497 863
rect 451 675 497 687
rect 609 863 655 875
rect 609 687 615 863
rect 649 687 655 863
rect 609 675 655 687
rect 767 863 813 875
rect 767 687 773 863
rect 807 687 813 863
rect 767 675 813 687
rect 925 863 971 875
rect 925 687 931 863
rect 965 687 971 863
rect 925 675 971 687
rect 1083 863 1129 875
rect 1083 687 1089 863
rect 1123 687 1129 863
rect 1083 675 1129 687
rect 1241 863 1287 875
rect 1241 687 1247 863
rect 1281 687 1287 863
rect 1241 675 1287 687
rect 1399 863 1445 875
rect 1399 687 1405 863
rect 1439 687 1445 863
rect 1399 675 1445 687
rect 1557 863 1603 875
rect 1557 687 1563 863
rect 1597 687 1603 863
rect 1557 675 1603 687
rect -1547 637 -1455 643
rect -1547 603 -1535 637
rect -1467 603 -1455 637
rect -1547 597 -1455 603
rect -1389 637 -1297 643
rect -1389 603 -1377 637
rect -1309 603 -1297 637
rect -1389 597 -1297 603
rect -1231 637 -1139 643
rect -1231 603 -1219 637
rect -1151 603 -1139 637
rect -1231 597 -1139 603
rect -1073 637 -981 643
rect -1073 603 -1061 637
rect -993 603 -981 637
rect -1073 597 -981 603
rect -915 637 -823 643
rect -915 603 -903 637
rect -835 603 -823 637
rect -915 597 -823 603
rect -757 637 -665 643
rect -757 603 -745 637
rect -677 603 -665 637
rect -757 597 -665 603
rect -599 637 -507 643
rect -599 603 -587 637
rect -519 603 -507 637
rect -599 597 -507 603
rect -441 637 -349 643
rect -441 603 -429 637
rect -361 603 -349 637
rect -441 597 -349 603
rect -283 637 -191 643
rect -283 603 -271 637
rect -203 603 -191 637
rect -283 597 -191 603
rect -125 637 -33 643
rect -125 603 -113 637
rect -45 603 -33 637
rect -125 597 -33 603
rect 33 637 125 643
rect 33 603 45 637
rect 113 603 125 637
rect 33 597 125 603
rect 191 637 283 643
rect 191 603 203 637
rect 271 603 283 637
rect 191 597 283 603
rect 349 637 441 643
rect 349 603 361 637
rect 429 603 441 637
rect 349 597 441 603
rect 507 637 599 643
rect 507 603 519 637
rect 587 603 599 637
rect 507 597 599 603
rect 665 637 757 643
rect 665 603 677 637
rect 745 603 757 637
rect 665 597 757 603
rect 823 637 915 643
rect 823 603 835 637
rect 903 603 915 637
rect 823 597 915 603
rect 981 637 1073 643
rect 981 603 993 637
rect 1061 603 1073 637
rect 981 597 1073 603
rect 1139 637 1231 643
rect 1139 603 1151 637
rect 1219 603 1231 637
rect 1139 597 1231 603
rect 1297 637 1389 643
rect 1297 603 1309 637
rect 1377 603 1389 637
rect 1297 597 1389 603
rect 1455 637 1547 643
rect 1455 603 1467 637
rect 1535 603 1547 637
rect 1455 597 1547 603
rect -1603 553 -1557 565
rect -1603 377 -1597 553
rect -1563 377 -1557 553
rect -1603 365 -1557 377
rect -1445 553 -1399 565
rect -1445 377 -1439 553
rect -1405 377 -1399 553
rect -1445 365 -1399 377
rect -1287 553 -1241 565
rect -1287 377 -1281 553
rect -1247 377 -1241 553
rect -1287 365 -1241 377
rect -1129 553 -1083 565
rect -1129 377 -1123 553
rect -1089 377 -1083 553
rect -1129 365 -1083 377
rect -971 553 -925 565
rect -971 377 -965 553
rect -931 377 -925 553
rect -971 365 -925 377
rect -813 553 -767 565
rect -813 377 -807 553
rect -773 377 -767 553
rect -813 365 -767 377
rect -655 553 -609 565
rect -655 377 -649 553
rect -615 377 -609 553
rect -655 365 -609 377
rect -497 553 -451 565
rect -497 377 -491 553
rect -457 377 -451 553
rect -497 365 -451 377
rect -339 553 -293 565
rect -339 377 -333 553
rect -299 377 -293 553
rect -339 365 -293 377
rect -181 553 -135 565
rect -181 377 -175 553
rect -141 377 -135 553
rect -181 365 -135 377
rect -23 553 23 565
rect -23 377 -17 553
rect 17 377 23 553
rect -23 365 23 377
rect 135 553 181 565
rect 135 377 141 553
rect 175 377 181 553
rect 135 365 181 377
rect 293 553 339 565
rect 293 377 299 553
rect 333 377 339 553
rect 293 365 339 377
rect 451 553 497 565
rect 451 377 457 553
rect 491 377 497 553
rect 451 365 497 377
rect 609 553 655 565
rect 609 377 615 553
rect 649 377 655 553
rect 609 365 655 377
rect 767 553 813 565
rect 767 377 773 553
rect 807 377 813 553
rect 767 365 813 377
rect 925 553 971 565
rect 925 377 931 553
rect 965 377 971 553
rect 925 365 971 377
rect 1083 553 1129 565
rect 1083 377 1089 553
rect 1123 377 1129 553
rect 1083 365 1129 377
rect 1241 553 1287 565
rect 1241 377 1247 553
rect 1281 377 1287 553
rect 1241 365 1287 377
rect 1399 553 1445 565
rect 1399 377 1405 553
rect 1439 377 1445 553
rect 1399 365 1445 377
rect 1557 553 1603 565
rect 1557 377 1563 553
rect 1597 377 1603 553
rect 1557 365 1603 377
rect -1547 327 -1455 333
rect -1547 293 -1535 327
rect -1467 293 -1455 327
rect -1547 287 -1455 293
rect -1389 327 -1297 333
rect -1389 293 -1377 327
rect -1309 293 -1297 327
rect -1389 287 -1297 293
rect -1231 327 -1139 333
rect -1231 293 -1219 327
rect -1151 293 -1139 327
rect -1231 287 -1139 293
rect -1073 327 -981 333
rect -1073 293 -1061 327
rect -993 293 -981 327
rect -1073 287 -981 293
rect -915 327 -823 333
rect -915 293 -903 327
rect -835 293 -823 327
rect -915 287 -823 293
rect -757 327 -665 333
rect -757 293 -745 327
rect -677 293 -665 327
rect -757 287 -665 293
rect -599 327 -507 333
rect -599 293 -587 327
rect -519 293 -507 327
rect -599 287 -507 293
rect -441 327 -349 333
rect -441 293 -429 327
rect -361 293 -349 327
rect -441 287 -349 293
rect -283 327 -191 333
rect -283 293 -271 327
rect -203 293 -191 327
rect -283 287 -191 293
rect -125 327 -33 333
rect -125 293 -113 327
rect -45 293 -33 327
rect -125 287 -33 293
rect 33 327 125 333
rect 33 293 45 327
rect 113 293 125 327
rect 33 287 125 293
rect 191 327 283 333
rect 191 293 203 327
rect 271 293 283 327
rect 191 287 283 293
rect 349 327 441 333
rect 349 293 361 327
rect 429 293 441 327
rect 349 287 441 293
rect 507 327 599 333
rect 507 293 519 327
rect 587 293 599 327
rect 507 287 599 293
rect 665 327 757 333
rect 665 293 677 327
rect 745 293 757 327
rect 665 287 757 293
rect 823 327 915 333
rect 823 293 835 327
rect 903 293 915 327
rect 823 287 915 293
rect 981 327 1073 333
rect 981 293 993 327
rect 1061 293 1073 327
rect 981 287 1073 293
rect 1139 327 1231 333
rect 1139 293 1151 327
rect 1219 293 1231 327
rect 1139 287 1231 293
rect 1297 327 1389 333
rect 1297 293 1309 327
rect 1377 293 1389 327
rect 1297 287 1389 293
rect 1455 327 1547 333
rect 1455 293 1467 327
rect 1535 293 1547 327
rect 1455 287 1547 293
rect -1603 243 -1557 255
rect -1603 67 -1597 243
rect -1563 67 -1557 243
rect -1603 55 -1557 67
rect -1445 243 -1399 255
rect -1445 67 -1439 243
rect -1405 67 -1399 243
rect -1445 55 -1399 67
rect -1287 243 -1241 255
rect -1287 67 -1281 243
rect -1247 67 -1241 243
rect -1287 55 -1241 67
rect -1129 243 -1083 255
rect -1129 67 -1123 243
rect -1089 67 -1083 243
rect -1129 55 -1083 67
rect -971 243 -925 255
rect -971 67 -965 243
rect -931 67 -925 243
rect -971 55 -925 67
rect -813 243 -767 255
rect -813 67 -807 243
rect -773 67 -767 243
rect -813 55 -767 67
rect -655 243 -609 255
rect -655 67 -649 243
rect -615 67 -609 243
rect -655 55 -609 67
rect -497 243 -451 255
rect -497 67 -491 243
rect -457 67 -451 243
rect -497 55 -451 67
rect -339 243 -293 255
rect -339 67 -333 243
rect -299 67 -293 243
rect -339 55 -293 67
rect -181 243 -135 255
rect -181 67 -175 243
rect -141 67 -135 243
rect -181 55 -135 67
rect -23 243 23 255
rect -23 67 -17 243
rect 17 67 23 243
rect -23 55 23 67
rect 135 243 181 255
rect 135 67 141 243
rect 175 67 181 243
rect 135 55 181 67
rect 293 243 339 255
rect 293 67 299 243
rect 333 67 339 243
rect 293 55 339 67
rect 451 243 497 255
rect 451 67 457 243
rect 491 67 497 243
rect 451 55 497 67
rect 609 243 655 255
rect 609 67 615 243
rect 649 67 655 243
rect 609 55 655 67
rect 767 243 813 255
rect 767 67 773 243
rect 807 67 813 243
rect 767 55 813 67
rect 925 243 971 255
rect 925 67 931 243
rect 965 67 971 243
rect 925 55 971 67
rect 1083 243 1129 255
rect 1083 67 1089 243
rect 1123 67 1129 243
rect 1083 55 1129 67
rect 1241 243 1287 255
rect 1241 67 1247 243
rect 1281 67 1287 243
rect 1241 55 1287 67
rect 1399 243 1445 255
rect 1399 67 1405 243
rect 1439 67 1445 243
rect 1399 55 1445 67
rect 1557 243 1603 255
rect 1557 67 1563 243
rect 1597 67 1603 243
rect 1557 55 1603 67
rect -1547 17 -1455 23
rect -1547 -17 -1535 17
rect -1467 -17 -1455 17
rect -1547 -23 -1455 -17
rect -1389 17 -1297 23
rect -1389 -17 -1377 17
rect -1309 -17 -1297 17
rect -1389 -23 -1297 -17
rect -1231 17 -1139 23
rect -1231 -17 -1219 17
rect -1151 -17 -1139 17
rect -1231 -23 -1139 -17
rect -1073 17 -981 23
rect -1073 -17 -1061 17
rect -993 -17 -981 17
rect -1073 -23 -981 -17
rect -915 17 -823 23
rect -915 -17 -903 17
rect -835 -17 -823 17
rect -915 -23 -823 -17
rect -757 17 -665 23
rect -757 -17 -745 17
rect -677 -17 -665 17
rect -757 -23 -665 -17
rect -599 17 -507 23
rect -599 -17 -587 17
rect -519 -17 -507 17
rect -599 -23 -507 -17
rect -441 17 -349 23
rect -441 -17 -429 17
rect -361 -17 -349 17
rect -441 -23 -349 -17
rect -283 17 -191 23
rect -283 -17 -271 17
rect -203 -17 -191 17
rect -283 -23 -191 -17
rect -125 17 -33 23
rect -125 -17 -113 17
rect -45 -17 -33 17
rect -125 -23 -33 -17
rect 33 17 125 23
rect 33 -17 45 17
rect 113 -17 125 17
rect 33 -23 125 -17
rect 191 17 283 23
rect 191 -17 203 17
rect 271 -17 283 17
rect 191 -23 283 -17
rect 349 17 441 23
rect 349 -17 361 17
rect 429 -17 441 17
rect 349 -23 441 -17
rect 507 17 599 23
rect 507 -17 519 17
rect 587 -17 599 17
rect 507 -23 599 -17
rect 665 17 757 23
rect 665 -17 677 17
rect 745 -17 757 17
rect 665 -23 757 -17
rect 823 17 915 23
rect 823 -17 835 17
rect 903 -17 915 17
rect 823 -23 915 -17
rect 981 17 1073 23
rect 981 -17 993 17
rect 1061 -17 1073 17
rect 981 -23 1073 -17
rect 1139 17 1231 23
rect 1139 -17 1151 17
rect 1219 -17 1231 17
rect 1139 -23 1231 -17
rect 1297 17 1389 23
rect 1297 -17 1309 17
rect 1377 -17 1389 17
rect 1297 -23 1389 -17
rect 1455 17 1547 23
rect 1455 -17 1467 17
rect 1535 -17 1547 17
rect 1455 -23 1547 -17
rect -1603 -67 -1557 -55
rect -1603 -243 -1597 -67
rect -1563 -243 -1557 -67
rect -1603 -255 -1557 -243
rect -1445 -67 -1399 -55
rect -1445 -243 -1439 -67
rect -1405 -243 -1399 -67
rect -1445 -255 -1399 -243
rect -1287 -67 -1241 -55
rect -1287 -243 -1281 -67
rect -1247 -243 -1241 -67
rect -1287 -255 -1241 -243
rect -1129 -67 -1083 -55
rect -1129 -243 -1123 -67
rect -1089 -243 -1083 -67
rect -1129 -255 -1083 -243
rect -971 -67 -925 -55
rect -971 -243 -965 -67
rect -931 -243 -925 -67
rect -971 -255 -925 -243
rect -813 -67 -767 -55
rect -813 -243 -807 -67
rect -773 -243 -767 -67
rect -813 -255 -767 -243
rect -655 -67 -609 -55
rect -655 -243 -649 -67
rect -615 -243 -609 -67
rect -655 -255 -609 -243
rect -497 -67 -451 -55
rect -497 -243 -491 -67
rect -457 -243 -451 -67
rect -497 -255 -451 -243
rect -339 -67 -293 -55
rect -339 -243 -333 -67
rect -299 -243 -293 -67
rect -339 -255 -293 -243
rect -181 -67 -135 -55
rect -181 -243 -175 -67
rect -141 -243 -135 -67
rect -181 -255 -135 -243
rect -23 -67 23 -55
rect -23 -243 -17 -67
rect 17 -243 23 -67
rect -23 -255 23 -243
rect 135 -67 181 -55
rect 135 -243 141 -67
rect 175 -243 181 -67
rect 135 -255 181 -243
rect 293 -67 339 -55
rect 293 -243 299 -67
rect 333 -243 339 -67
rect 293 -255 339 -243
rect 451 -67 497 -55
rect 451 -243 457 -67
rect 491 -243 497 -67
rect 451 -255 497 -243
rect 609 -67 655 -55
rect 609 -243 615 -67
rect 649 -243 655 -67
rect 609 -255 655 -243
rect 767 -67 813 -55
rect 767 -243 773 -67
rect 807 -243 813 -67
rect 767 -255 813 -243
rect 925 -67 971 -55
rect 925 -243 931 -67
rect 965 -243 971 -67
rect 925 -255 971 -243
rect 1083 -67 1129 -55
rect 1083 -243 1089 -67
rect 1123 -243 1129 -67
rect 1083 -255 1129 -243
rect 1241 -67 1287 -55
rect 1241 -243 1247 -67
rect 1281 -243 1287 -67
rect 1241 -255 1287 -243
rect 1399 -67 1445 -55
rect 1399 -243 1405 -67
rect 1439 -243 1445 -67
rect 1399 -255 1445 -243
rect 1557 -67 1603 -55
rect 1557 -243 1563 -67
rect 1597 -243 1603 -67
rect 1557 -255 1603 -243
rect -1547 -293 -1455 -287
rect -1547 -327 -1535 -293
rect -1467 -327 -1455 -293
rect -1547 -333 -1455 -327
rect -1389 -293 -1297 -287
rect -1389 -327 -1377 -293
rect -1309 -327 -1297 -293
rect -1389 -333 -1297 -327
rect -1231 -293 -1139 -287
rect -1231 -327 -1219 -293
rect -1151 -327 -1139 -293
rect -1231 -333 -1139 -327
rect -1073 -293 -981 -287
rect -1073 -327 -1061 -293
rect -993 -327 -981 -293
rect -1073 -333 -981 -327
rect -915 -293 -823 -287
rect -915 -327 -903 -293
rect -835 -327 -823 -293
rect -915 -333 -823 -327
rect -757 -293 -665 -287
rect -757 -327 -745 -293
rect -677 -327 -665 -293
rect -757 -333 -665 -327
rect -599 -293 -507 -287
rect -599 -327 -587 -293
rect -519 -327 -507 -293
rect -599 -333 -507 -327
rect -441 -293 -349 -287
rect -441 -327 -429 -293
rect -361 -327 -349 -293
rect -441 -333 -349 -327
rect -283 -293 -191 -287
rect -283 -327 -271 -293
rect -203 -327 -191 -293
rect -283 -333 -191 -327
rect -125 -293 -33 -287
rect -125 -327 -113 -293
rect -45 -327 -33 -293
rect -125 -333 -33 -327
rect 33 -293 125 -287
rect 33 -327 45 -293
rect 113 -327 125 -293
rect 33 -333 125 -327
rect 191 -293 283 -287
rect 191 -327 203 -293
rect 271 -327 283 -293
rect 191 -333 283 -327
rect 349 -293 441 -287
rect 349 -327 361 -293
rect 429 -327 441 -293
rect 349 -333 441 -327
rect 507 -293 599 -287
rect 507 -327 519 -293
rect 587 -327 599 -293
rect 507 -333 599 -327
rect 665 -293 757 -287
rect 665 -327 677 -293
rect 745 -327 757 -293
rect 665 -333 757 -327
rect 823 -293 915 -287
rect 823 -327 835 -293
rect 903 -327 915 -293
rect 823 -333 915 -327
rect 981 -293 1073 -287
rect 981 -327 993 -293
rect 1061 -327 1073 -293
rect 981 -333 1073 -327
rect 1139 -293 1231 -287
rect 1139 -327 1151 -293
rect 1219 -327 1231 -293
rect 1139 -333 1231 -327
rect 1297 -293 1389 -287
rect 1297 -327 1309 -293
rect 1377 -327 1389 -293
rect 1297 -333 1389 -327
rect 1455 -293 1547 -287
rect 1455 -327 1467 -293
rect 1535 -327 1547 -293
rect 1455 -333 1547 -327
rect -1603 -377 -1557 -365
rect -1603 -553 -1597 -377
rect -1563 -553 -1557 -377
rect -1603 -565 -1557 -553
rect -1445 -377 -1399 -365
rect -1445 -553 -1439 -377
rect -1405 -553 -1399 -377
rect -1445 -565 -1399 -553
rect -1287 -377 -1241 -365
rect -1287 -553 -1281 -377
rect -1247 -553 -1241 -377
rect -1287 -565 -1241 -553
rect -1129 -377 -1083 -365
rect -1129 -553 -1123 -377
rect -1089 -553 -1083 -377
rect -1129 -565 -1083 -553
rect -971 -377 -925 -365
rect -971 -553 -965 -377
rect -931 -553 -925 -377
rect -971 -565 -925 -553
rect -813 -377 -767 -365
rect -813 -553 -807 -377
rect -773 -553 -767 -377
rect -813 -565 -767 -553
rect -655 -377 -609 -365
rect -655 -553 -649 -377
rect -615 -553 -609 -377
rect -655 -565 -609 -553
rect -497 -377 -451 -365
rect -497 -553 -491 -377
rect -457 -553 -451 -377
rect -497 -565 -451 -553
rect -339 -377 -293 -365
rect -339 -553 -333 -377
rect -299 -553 -293 -377
rect -339 -565 -293 -553
rect -181 -377 -135 -365
rect -181 -553 -175 -377
rect -141 -553 -135 -377
rect -181 -565 -135 -553
rect -23 -377 23 -365
rect -23 -553 -17 -377
rect 17 -553 23 -377
rect -23 -565 23 -553
rect 135 -377 181 -365
rect 135 -553 141 -377
rect 175 -553 181 -377
rect 135 -565 181 -553
rect 293 -377 339 -365
rect 293 -553 299 -377
rect 333 -553 339 -377
rect 293 -565 339 -553
rect 451 -377 497 -365
rect 451 -553 457 -377
rect 491 -553 497 -377
rect 451 -565 497 -553
rect 609 -377 655 -365
rect 609 -553 615 -377
rect 649 -553 655 -377
rect 609 -565 655 -553
rect 767 -377 813 -365
rect 767 -553 773 -377
rect 807 -553 813 -377
rect 767 -565 813 -553
rect 925 -377 971 -365
rect 925 -553 931 -377
rect 965 -553 971 -377
rect 925 -565 971 -553
rect 1083 -377 1129 -365
rect 1083 -553 1089 -377
rect 1123 -553 1129 -377
rect 1083 -565 1129 -553
rect 1241 -377 1287 -365
rect 1241 -553 1247 -377
rect 1281 -553 1287 -377
rect 1241 -565 1287 -553
rect 1399 -377 1445 -365
rect 1399 -553 1405 -377
rect 1439 -553 1445 -377
rect 1399 -565 1445 -553
rect 1557 -377 1603 -365
rect 1557 -553 1563 -377
rect 1597 -553 1603 -377
rect 1557 -565 1603 -553
rect -1547 -603 -1455 -597
rect -1547 -637 -1535 -603
rect -1467 -637 -1455 -603
rect -1547 -643 -1455 -637
rect -1389 -603 -1297 -597
rect -1389 -637 -1377 -603
rect -1309 -637 -1297 -603
rect -1389 -643 -1297 -637
rect -1231 -603 -1139 -597
rect -1231 -637 -1219 -603
rect -1151 -637 -1139 -603
rect -1231 -643 -1139 -637
rect -1073 -603 -981 -597
rect -1073 -637 -1061 -603
rect -993 -637 -981 -603
rect -1073 -643 -981 -637
rect -915 -603 -823 -597
rect -915 -637 -903 -603
rect -835 -637 -823 -603
rect -915 -643 -823 -637
rect -757 -603 -665 -597
rect -757 -637 -745 -603
rect -677 -637 -665 -603
rect -757 -643 -665 -637
rect -599 -603 -507 -597
rect -599 -637 -587 -603
rect -519 -637 -507 -603
rect -599 -643 -507 -637
rect -441 -603 -349 -597
rect -441 -637 -429 -603
rect -361 -637 -349 -603
rect -441 -643 -349 -637
rect -283 -603 -191 -597
rect -283 -637 -271 -603
rect -203 -637 -191 -603
rect -283 -643 -191 -637
rect -125 -603 -33 -597
rect -125 -637 -113 -603
rect -45 -637 -33 -603
rect -125 -643 -33 -637
rect 33 -603 125 -597
rect 33 -637 45 -603
rect 113 -637 125 -603
rect 33 -643 125 -637
rect 191 -603 283 -597
rect 191 -637 203 -603
rect 271 -637 283 -603
rect 191 -643 283 -637
rect 349 -603 441 -597
rect 349 -637 361 -603
rect 429 -637 441 -603
rect 349 -643 441 -637
rect 507 -603 599 -597
rect 507 -637 519 -603
rect 587 -637 599 -603
rect 507 -643 599 -637
rect 665 -603 757 -597
rect 665 -637 677 -603
rect 745 -637 757 -603
rect 665 -643 757 -637
rect 823 -603 915 -597
rect 823 -637 835 -603
rect 903 -637 915 -603
rect 823 -643 915 -637
rect 981 -603 1073 -597
rect 981 -637 993 -603
rect 1061 -637 1073 -603
rect 981 -643 1073 -637
rect 1139 -603 1231 -597
rect 1139 -637 1151 -603
rect 1219 -637 1231 -603
rect 1139 -643 1231 -637
rect 1297 -603 1389 -597
rect 1297 -637 1309 -603
rect 1377 -637 1389 -603
rect 1297 -643 1389 -637
rect 1455 -603 1547 -597
rect 1455 -637 1467 -603
rect 1535 -637 1547 -603
rect 1455 -643 1547 -637
rect -1603 -687 -1557 -675
rect -1603 -863 -1597 -687
rect -1563 -863 -1557 -687
rect -1603 -875 -1557 -863
rect -1445 -687 -1399 -675
rect -1445 -863 -1439 -687
rect -1405 -863 -1399 -687
rect -1445 -875 -1399 -863
rect -1287 -687 -1241 -675
rect -1287 -863 -1281 -687
rect -1247 -863 -1241 -687
rect -1287 -875 -1241 -863
rect -1129 -687 -1083 -675
rect -1129 -863 -1123 -687
rect -1089 -863 -1083 -687
rect -1129 -875 -1083 -863
rect -971 -687 -925 -675
rect -971 -863 -965 -687
rect -931 -863 -925 -687
rect -971 -875 -925 -863
rect -813 -687 -767 -675
rect -813 -863 -807 -687
rect -773 -863 -767 -687
rect -813 -875 -767 -863
rect -655 -687 -609 -675
rect -655 -863 -649 -687
rect -615 -863 -609 -687
rect -655 -875 -609 -863
rect -497 -687 -451 -675
rect -497 -863 -491 -687
rect -457 -863 -451 -687
rect -497 -875 -451 -863
rect -339 -687 -293 -675
rect -339 -863 -333 -687
rect -299 -863 -293 -687
rect -339 -875 -293 -863
rect -181 -687 -135 -675
rect -181 -863 -175 -687
rect -141 -863 -135 -687
rect -181 -875 -135 -863
rect -23 -687 23 -675
rect -23 -863 -17 -687
rect 17 -863 23 -687
rect -23 -875 23 -863
rect 135 -687 181 -675
rect 135 -863 141 -687
rect 175 -863 181 -687
rect 135 -875 181 -863
rect 293 -687 339 -675
rect 293 -863 299 -687
rect 333 -863 339 -687
rect 293 -875 339 -863
rect 451 -687 497 -675
rect 451 -863 457 -687
rect 491 -863 497 -687
rect 451 -875 497 -863
rect 609 -687 655 -675
rect 609 -863 615 -687
rect 649 -863 655 -687
rect 609 -875 655 -863
rect 767 -687 813 -675
rect 767 -863 773 -687
rect 807 -863 813 -687
rect 767 -875 813 -863
rect 925 -687 971 -675
rect 925 -863 931 -687
rect 965 -863 971 -687
rect 925 -875 971 -863
rect 1083 -687 1129 -675
rect 1083 -863 1089 -687
rect 1123 -863 1129 -687
rect 1083 -875 1129 -863
rect 1241 -687 1287 -675
rect 1241 -863 1247 -687
rect 1281 -863 1287 -687
rect 1241 -875 1287 -863
rect 1399 -687 1445 -675
rect 1399 -863 1405 -687
rect 1439 -863 1445 -687
rect 1399 -875 1445 -863
rect 1557 -687 1603 -675
rect 1557 -863 1563 -687
rect 1597 -863 1603 -687
rect 1557 -875 1603 -863
rect -1547 -913 -1455 -907
rect -1547 -947 -1535 -913
rect -1467 -947 -1455 -913
rect -1547 -953 -1455 -947
rect -1389 -913 -1297 -907
rect -1389 -947 -1377 -913
rect -1309 -947 -1297 -913
rect -1389 -953 -1297 -947
rect -1231 -913 -1139 -907
rect -1231 -947 -1219 -913
rect -1151 -947 -1139 -913
rect -1231 -953 -1139 -947
rect -1073 -913 -981 -907
rect -1073 -947 -1061 -913
rect -993 -947 -981 -913
rect -1073 -953 -981 -947
rect -915 -913 -823 -907
rect -915 -947 -903 -913
rect -835 -947 -823 -913
rect -915 -953 -823 -947
rect -757 -913 -665 -907
rect -757 -947 -745 -913
rect -677 -947 -665 -913
rect -757 -953 -665 -947
rect -599 -913 -507 -907
rect -599 -947 -587 -913
rect -519 -947 -507 -913
rect -599 -953 -507 -947
rect -441 -913 -349 -907
rect -441 -947 -429 -913
rect -361 -947 -349 -913
rect -441 -953 -349 -947
rect -283 -913 -191 -907
rect -283 -947 -271 -913
rect -203 -947 -191 -913
rect -283 -953 -191 -947
rect -125 -913 -33 -907
rect -125 -947 -113 -913
rect -45 -947 -33 -913
rect -125 -953 -33 -947
rect 33 -913 125 -907
rect 33 -947 45 -913
rect 113 -947 125 -913
rect 33 -953 125 -947
rect 191 -913 283 -907
rect 191 -947 203 -913
rect 271 -947 283 -913
rect 191 -953 283 -947
rect 349 -913 441 -907
rect 349 -947 361 -913
rect 429 -947 441 -913
rect 349 -953 441 -947
rect 507 -913 599 -907
rect 507 -947 519 -913
rect 587 -947 599 -913
rect 507 -953 599 -947
rect 665 -913 757 -907
rect 665 -947 677 -913
rect 745 -947 757 -913
rect 665 -953 757 -947
rect 823 -913 915 -907
rect 823 -947 835 -913
rect 903 -947 915 -913
rect 823 -953 915 -947
rect 981 -913 1073 -907
rect 981 -947 993 -913
rect 1061 -947 1073 -913
rect 981 -953 1073 -947
rect 1139 -913 1231 -907
rect 1139 -947 1151 -913
rect 1219 -947 1231 -913
rect 1139 -953 1231 -947
rect 1297 -913 1389 -907
rect 1297 -947 1309 -913
rect 1377 -947 1389 -913
rect 1297 -953 1389 -947
rect 1455 -913 1547 -907
rect 1455 -947 1467 -913
rect 1535 -947 1547 -913
rect 1455 -953 1547 -947
rect -1603 -997 -1557 -985
rect -1603 -1173 -1597 -997
rect -1563 -1173 -1557 -997
rect -1603 -1185 -1557 -1173
rect -1445 -997 -1399 -985
rect -1445 -1173 -1439 -997
rect -1405 -1173 -1399 -997
rect -1445 -1185 -1399 -1173
rect -1287 -997 -1241 -985
rect -1287 -1173 -1281 -997
rect -1247 -1173 -1241 -997
rect -1287 -1185 -1241 -1173
rect -1129 -997 -1083 -985
rect -1129 -1173 -1123 -997
rect -1089 -1173 -1083 -997
rect -1129 -1185 -1083 -1173
rect -971 -997 -925 -985
rect -971 -1173 -965 -997
rect -931 -1173 -925 -997
rect -971 -1185 -925 -1173
rect -813 -997 -767 -985
rect -813 -1173 -807 -997
rect -773 -1173 -767 -997
rect -813 -1185 -767 -1173
rect -655 -997 -609 -985
rect -655 -1173 -649 -997
rect -615 -1173 -609 -997
rect -655 -1185 -609 -1173
rect -497 -997 -451 -985
rect -497 -1173 -491 -997
rect -457 -1173 -451 -997
rect -497 -1185 -451 -1173
rect -339 -997 -293 -985
rect -339 -1173 -333 -997
rect -299 -1173 -293 -997
rect -339 -1185 -293 -1173
rect -181 -997 -135 -985
rect -181 -1173 -175 -997
rect -141 -1173 -135 -997
rect -181 -1185 -135 -1173
rect -23 -997 23 -985
rect -23 -1173 -17 -997
rect 17 -1173 23 -997
rect -23 -1185 23 -1173
rect 135 -997 181 -985
rect 135 -1173 141 -997
rect 175 -1173 181 -997
rect 135 -1185 181 -1173
rect 293 -997 339 -985
rect 293 -1173 299 -997
rect 333 -1173 339 -997
rect 293 -1185 339 -1173
rect 451 -997 497 -985
rect 451 -1173 457 -997
rect 491 -1173 497 -997
rect 451 -1185 497 -1173
rect 609 -997 655 -985
rect 609 -1173 615 -997
rect 649 -1173 655 -997
rect 609 -1185 655 -1173
rect 767 -997 813 -985
rect 767 -1173 773 -997
rect 807 -1173 813 -997
rect 767 -1185 813 -1173
rect 925 -997 971 -985
rect 925 -1173 931 -997
rect 965 -1173 971 -997
rect 925 -1185 971 -1173
rect 1083 -997 1129 -985
rect 1083 -1173 1089 -997
rect 1123 -1173 1129 -997
rect 1083 -1185 1129 -1173
rect 1241 -997 1287 -985
rect 1241 -1173 1247 -997
rect 1281 -1173 1287 -997
rect 1241 -1185 1287 -1173
rect 1399 -997 1445 -985
rect 1399 -1173 1405 -997
rect 1439 -1173 1445 -997
rect 1399 -1185 1445 -1173
rect 1557 -997 1603 -985
rect 1557 -1173 1563 -997
rect 1597 -1173 1603 -997
rect 1557 -1185 1603 -1173
rect -1547 -1223 -1455 -1217
rect -1547 -1257 -1535 -1223
rect -1467 -1257 -1455 -1223
rect -1547 -1263 -1455 -1257
rect -1389 -1223 -1297 -1217
rect -1389 -1257 -1377 -1223
rect -1309 -1257 -1297 -1223
rect -1389 -1263 -1297 -1257
rect -1231 -1223 -1139 -1217
rect -1231 -1257 -1219 -1223
rect -1151 -1257 -1139 -1223
rect -1231 -1263 -1139 -1257
rect -1073 -1223 -981 -1217
rect -1073 -1257 -1061 -1223
rect -993 -1257 -981 -1223
rect -1073 -1263 -981 -1257
rect -915 -1223 -823 -1217
rect -915 -1257 -903 -1223
rect -835 -1257 -823 -1223
rect -915 -1263 -823 -1257
rect -757 -1223 -665 -1217
rect -757 -1257 -745 -1223
rect -677 -1257 -665 -1223
rect -757 -1263 -665 -1257
rect -599 -1223 -507 -1217
rect -599 -1257 -587 -1223
rect -519 -1257 -507 -1223
rect -599 -1263 -507 -1257
rect -441 -1223 -349 -1217
rect -441 -1257 -429 -1223
rect -361 -1257 -349 -1223
rect -441 -1263 -349 -1257
rect -283 -1223 -191 -1217
rect -283 -1257 -271 -1223
rect -203 -1257 -191 -1223
rect -283 -1263 -191 -1257
rect -125 -1223 -33 -1217
rect -125 -1257 -113 -1223
rect -45 -1257 -33 -1223
rect -125 -1263 -33 -1257
rect 33 -1223 125 -1217
rect 33 -1257 45 -1223
rect 113 -1257 125 -1223
rect 33 -1263 125 -1257
rect 191 -1223 283 -1217
rect 191 -1257 203 -1223
rect 271 -1257 283 -1223
rect 191 -1263 283 -1257
rect 349 -1223 441 -1217
rect 349 -1257 361 -1223
rect 429 -1257 441 -1223
rect 349 -1263 441 -1257
rect 507 -1223 599 -1217
rect 507 -1257 519 -1223
rect 587 -1257 599 -1223
rect 507 -1263 599 -1257
rect 665 -1223 757 -1217
rect 665 -1257 677 -1223
rect 745 -1257 757 -1223
rect 665 -1263 757 -1257
rect 823 -1223 915 -1217
rect 823 -1257 835 -1223
rect 903 -1257 915 -1223
rect 823 -1263 915 -1257
rect 981 -1223 1073 -1217
rect 981 -1257 993 -1223
rect 1061 -1257 1073 -1223
rect 981 -1263 1073 -1257
rect 1139 -1223 1231 -1217
rect 1139 -1257 1151 -1223
rect 1219 -1257 1231 -1223
rect 1139 -1263 1231 -1257
rect 1297 -1223 1389 -1217
rect 1297 -1257 1309 -1223
rect 1377 -1257 1389 -1223
rect 1297 -1263 1389 -1257
rect 1455 -1223 1547 -1217
rect 1455 -1257 1467 -1223
rect 1535 -1257 1547 -1223
rect 1455 -1263 1547 -1257
rect -1603 -1307 -1557 -1295
rect -1603 -1483 -1597 -1307
rect -1563 -1483 -1557 -1307
rect -1603 -1495 -1557 -1483
rect -1445 -1307 -1399 -1295
rect -1445 -1483 -1439 -1307
rect -1405 -1483 -1399 -1307
rect -1445 -1495 -1399 -1483
rect -1287 -1307 -1241 -1295
rect -1287 -1483 -1281 -1307
rect -1247 -1483 -1241 -1307
rect -1287 -1495 -1241 -1483
rect -1129 -1307 -1083 -1295
rect -1129 -1483 -1123 -1307
rect -1089 -1483 -1083 -1307
rect -1129 -1495 -1083 -1483
rect -971 -1307 -925 -1295
rect -971 -1483 -965 -1307
rect -931 -1483 -925 -1307
rect -971 -1495 -925 -1483
rect -813 -1307 -767 -1295
rect -813 -1483 -807 -1307
rect -773 -1483 -767 -1307
rect -813 -1495 -767 -1483
rect -655 -1307 -609 -1295
rect -655 -1483 -649 -1307
rect -615 -1483 -609 -1307
rect -655 -1495 -609 -1483
rect -497 -1307 -451 -1295
rect -497 -1483 -491 -1307
rect -457 -1483 -451 -1307
rect -497 -1495 -451 -1483
rect -339 -1307 -293 -1295
rect -339 -1483 -333 -1307
rect -299 -1483 -293 -1307
rect -339 -1495 -293 -1483
rect -181 -1307 -135 -1295
rect -181 -1483 -175 -1307
rect -141 -1483 -135 -1307
rect -181 -1495 -135 -1483
rect -23 -1307 23 -1295
rect -23 -1483 -17 -1307
rect 17 -1483 23 -1307
rect -23 -1495 23 -1483
rect 135 -1307 181 -1295
rect 135 -1483 141 -1307
rect 175 -1483 181 -1307
rect 135 -1495 181 -1483
rect 293 -1307 339 -1295
rect 293 -1483 299 -1307
rect 333 -1483 339 -1307
rect 293 -1495 339 -1483
rect 451 -1307 497 -1295
rect 451 -1483 457 -1307
rect 491 -1483 497 -1307
rect 451 -1495 497 -1483
rect 609 -1307 655 -1295
rect 609 -1483 615 -1307
rect 649 -1483 655 -1307
rect 609 -1495 655 -1483
rect 767 -1307 813 -1295
rect 767 -1483 773 -1307
rect 807 -1483 813 -1307
rect 767 -1495 813 -1483
rect 925 -1307 971 -1295
rect 925 -1483 931 -1307
rect 965 -1483 971 -1307
rect 925 -1495 971 -1483
rect 1083 -1307 1129 -1295
rect 1083 -1483 1089 -1307
rect 1123 -1483 1129 -1307
rect 1083 -1495 1129 -1483
rect 1241 -1307 1287 -1295
rect 1241 -1483 1247 -1307
rect 1281 -1483 1287 -1307
rect 1241 -1495 1287 -1483
rect 1399 -1307 1445 -1295
rect 1399 -1483 1405 -1307
rect 1439 -1483 1445 -1307
rect 1399 -1495 1445 -1483
rect 1557 -1307 1603 -1295
rect 1557 -1483 1563 -1307
rect 1597 -1483 1603 -1307
rect 1557 -1495 1603 -1483
rect -1547 -1533 -1455 -1527
rect -1547 -1567 -1535 -1533
rect -1467 -1567 -1455 -1533
rect -1547 -1573 -1455 -1567
rect -1389 -1533 -1297 -1527
rect -1389 -1567 -1377 -1533
rect -1309 -1567 -1297 -1533
rect -1389 -1573 -1297 -1567
rect -1231 -1533 -1139 -1527
rect -1231 -1567 -1219 -1533
rect -1151 -1567 -1139 -1533
rect -1231 -1573 -1139 -1567
rect -1073 -1533 -981 -1527
rect -1073 -1567 -1061 -1533
rect -993 -1567 -981 -1533
rect -1073 -1573 -981 -1567
rect -915 -1533 -823 -1527
rect -915 -1567 -903 -1533
rect -835 -1567 -823 -1533
rect -915 -1573 -823 -1567
rect -757 -1533 -665 -1527
rect -757 -1567 -745 -1533
rect -677 -1567 -665 -1533
rect -757 -1573 -665 -1567
rect -599 -1533 -507 -1527
rect -599 -1567 -587 -1533
rect -519 -1567 -507 -1533
rect -599 -1573 -507 -1567
rect -441 -1533 -349 -1527
rect -441 -1567 -429 -1533
rect -361 -1567 -349 -1533
rect -441 -1573 -349 -1567
rect -283 -1533 -191 -1527
rect -283 -1567 -271 -1533
rect -203 -1567 -191 -1533
rect -283 -1573 -191 -1567
rect -125 -1533 -33 -1527
rect -125 -1567 -113 -1533
rect -45 -1567 -33 -1533
rect -125 -1573 -33 -1567
rect 33 -1533 125 -1527
rect 33 -1567 45 -1533
rect 113 -1567 125 -1533
rect 33 -1573 125 -1567
rect 191 -1533 283 -1527
rect 191 -1567 203 -1533
rect 271 -1567 283 -1533
rect 191 -1573 283 -1567
rect 349 -1533 441 -1527
rect 349 -1567 361 -1533
rect 429 -1567 441 -1533
rect 349 -1573 441 -1567
rect 507 -1533 599 -1527
rect 507 -1567 519 -1533
rect 587 -1567 599 -1533
rect 507 -1573 599 -1567
rect 665 -1533 757 -1527
rect 665 -1567 677 -1533
rect 745 -1567 757 -1533
rect 665 -1573 757 -1567
rect 823 -1533 915 -1527
rect 823 -1567 835 -1533
rect 903 -1567 915 -1533
rect 823 -1573 915 -1567
rect 981 -1533 1073 -1527
rect 981 -1567 993 -1533
rect 1061 -1567 1073 -1533
rect 981 -1573 1073 -1567
rect 1139 -1533 1231 -1527
rect 1139 -1567 1151 -1533
rect 1219 -1567 1231 -1533
rect 1139 -1573 1231 -1567
rect 1297 -1533 1389 -1527
rect 1297 -1567 1309 -1533
rect 1377 -1567 1389 -1533
rect 1297 -1573 1389 -1567
rect 1455 -1533 1547 -1527
rect 1455 -1567 1467 -1533
rect 1535 -1567 1547 -1533
rect 1455 -1573 1547 -1567
<< properties >>
string FIXED_BBOX -1714 -1688 1714 1688
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.50 m 10 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
