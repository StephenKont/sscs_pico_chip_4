magic
tech sky130A
magscale 1 2
timestamp 1666808413
<< viali >>
rect 1954 19740 1990 19782
rect 1956 19076 1992 19118
rect 1954 18966 1990 19008
rect 1954 18884 1990 18926
rect 1954 18288 1990 18330
rect 1954 18102 1990 18144
rect 1956 17446 1992 17488
rect 1956 17278 1992 17320
rect 1954 16586 1990 16628
rect 1954 16394 1990 16436
rect 1956 15778 1992 15820
rect 1954 15690 1990 15732
rect 1956 15542 1992 15584
rect 1956 14928 1992 14970
rect 1954 14830 1990 14872
rect 1954 14736 1990 14778
rect 1954 14644 1990 14686
rect 1956 13994 1992 14036
rect 1954 13834 1990 13876
rect 1954 13742 1990 13784
rect 1954 13134 1990 13176
rect 1954 13034 1990 13076
rect 1954 12356 1990 12398
rect 1956 12224 1992 12266
rect 1954 12108 1990 12150
rect 1956 11946 1992 11988
<< metal1 >>
rect 2118 19948 14048 20058
rect 2036 19808 2146 19898
rect 1940 19782 2146 19808
rect 1940 19740 1954 19782
rect 1990 19740 2146 19782
rect 1940 19720 2146 19740
rect 1942 19664 2146 19720
rect 1942 19184 2084 19664
rect 2140 19184 2146 19664
rect 1942 19118 2146 19184
rect 1942 19076 1956 19118
rect 1992 19076 2146 19118
rect 1942 19008 2146 19076
rect 1942 18966 1954 19008
rect 1990 18966 2146 19008
rect 1942 18926 2146 18966
rect 1942 18884 1954 18926
rect 1990 18884 2146 18926
rect 1942 18330 2146 18884
rect 1942 18288 1954 18330
rect 1990 18288 2146 18330
rect 1942 18144 2146 18288
rect 1942 18102 1954 18144
rect 1990 18102 2146 18144
rect 1942 18048 2146 18102
rect 1942 17568 2072 18048
rect 2128 17568 2146 18048
rect 1942 17488 2146 17568
rect 1942 17446 1956 17488
rect 1992 17446 2146 17488
rect 1942 17320 2146 17446
rect 1942 17278 1956 17320
rect 1992 17278 2146 17320
rect 1942 16628 2146 17278
rect 1942 16586 1954 16628
rect 1990 16586 2146 16628
rect 1942 16436 2146 16586
rect 1942 16394 1954 16436
rect 1990 16394 2146 16436
rect 1942 16326 2146 16394
rect 1942 15846 2066 16326
rect 2122 15846 2146 16326
rect 1942 15820 2146 15846
rect 1942 15778 1956 15820
rect 1992 15778 2146 15820
rect 1942 15732 2146 15778
rect 1942 15690 1954 15732
rect 1990 15690 2146 15732
rect 1942 15584 2146 15690
rect 1942 15542 1956 15584
rect 1992 15542 2146 15584
rect 1942 14970 2146 15542
rect 1942 14928 1956 14970
rect 1992 14928 2146 14970
rect 1942 14872 2146 14928
rect 1942 14830 1954 14872
rect 1990 14830 2146 14872
rect 1942 14778 2146 14830
rect 1942 14736 1954 14778
rect 1990 14736 2146 14778
rect 1942 14686 2146 14736
rect 1942 14644 1954 14686
rect 1990 14644 2146 14686
rect 1942 14544 2146 14644
rect 1942 14064 2076 14544
rect 2132 14064 2146 14544
rect 1942 14036 2146 14064
rect 1942 13994 1956 14036
rect 1992 13994 2146 14036
rect 1942 13876 2146 13994
rect 1942 13834 1954 13876
rect 1990 13834 2146 13876
rect 1942 13784 2146 13834
rect 1942 13742 1954 13784
rect 1990 13742 2146 13784
rect 1942 13176 2146 13742
rect 1942 13134 1954 13176
rect 1990 13134 2146 13176
rect 1942 13076 2146 13134
rect 1942 13034 1954 13076
rect 1990 13034 2146 13076
rect 1942 12928 2146 13034
rect 1942 12448 2066 12928
rect 2122 12448 2146 12928
rect 1942 12398 2146 12448
rect 1942 12356 1954 12398
rect 1990 12356 2146 12398
rect 1942 12266 2146 12356
rect 1942 12224 1956 12266
rect 1992 12224 2146 12266
rect 1942 12150 2146 12224
rect 1942 12108 1954 12150
rect 1990 12108 2146 12150
rect 1942 11988 2146 12108
rect 1942 11946 1956 11988
rect 1992 11946 2146 11988
rect 1942 11906 2146 11946
rect 2036 11898 2146 11906
rect 2222 18846 2316 19888
rect 2222 18366 2234 18846
rect 2290 18366 2316 18846
rect 2222 17208 2316 18366
rect 2222 16728 2236 17208
rect 2292 16728 2316 17208
rect 2222 15488 2316 16728
rect 2222 15008 2234 15488
rect 2290 15008 2316 15488
rect 2222 13692 2316 15008
rect 2222 13212 2226 13692
rect 2282 13212 2316 13692
rect 2222 11902 2316 13212
rect 2680 19676 2750 19884
rect 2680 19664 2760 19676
rect 2680 19184 2694 19664
rect 2750 19184 2760 19664
rect 2680 19174 2760 19184
rect 2680 18060 2750 19174
rect 2842 18858 2936 19888
rect 3298 19676 3368 19872
rect 3294 19664 3370 19676
rect 3294 19184 3304 19664
rect 3360 19184 3370 19664
rect 3294 19174 3370 19184
rect 2816 18844 2936 18858
rect 2816 18364 2852 18844
rect 2908 18364 2936 18844
rect 2816 18358 2936 18364
rect 2680 17580 2688 18060
rect 2744 17580 2750 18060
rect 2680 16322 2750 17580
rect 2680 15842 2688 16322
rect 2744 15842 2750 16322
rect 2680 14548 2750 15842
rect 2680 14068 2688 14548
rect 2744 14068 2750 14548
rect 2680 12918 2750 14068
rect 2680 12438 2688 12918
rect 2744 12438 2750 12918
rect 2680 11908 2750 12438
rect 2842 17194 2936 18358
rect 2842 16714 2852 17194
rect 2908 16714 2936 17194
rect 2842 15474 2936 16714
rect 2842 14994 2854 15474
rect 2910 14994 2936 15474
rect 2842 13686 2936 14994
rect 2842 13206 2848 13686
rect 2904 13206 2936 13686
rect 2842 11902 2936 13206
rect 3298 18060 3368 19174
rect 3460 18864 3536 19902
rect 3912 19676 3982 19876
rect 3912 19664 4000 19676
rect 3912 19184 3924 19664
rect 3980 19184 4000 19664
rect 3912 19176 4000 19184
rect 3458 18852 3560 18864
rect 3458 18372 3470 18852
rect 3526 18372 3560 18852
rect 3458 18364 3560 18372
rect 3460 18358 3556 18364
rect 3298 17580 3308 18060
rect 3364 17580 3368 18060
rect 3298 16326 3368 17580
rect 3298 15846 3312 16326
rect 3298 14544 3368 15846
rect 3298 14064 3308 14544
rect 3364 14064 3368 14544
rect 3298 12926 3368 14064
rect 3298 12446 3308 12926
rect 3364 12446 3368 12926
rect 3298 11896 3368 12446
rect 3462 17210 3556 18358
rect 3462 16730 3478 17210
rect 3534 16730 3556 17210
rect 3462 15488 3556 16730
rect 3462 15008 3474 15488
rect 3530 15008 3556 15488
rect 3462 13700 3556 15008
rect 3462 13220 3470 13700
rect 3526 13220 3556 13700
rect 3462 11902 3556 13220
rect 3912 18060 3982 19176
rect 4072 18842 4158 19898
rect 4530 19676 4600 19878
rect 4526 19664 4610 19676
rect 4526 19184 4534 19664
rect 4600 19184 4610 19664
rect 4526 19176 4610 19184
rect 4072 18362 4084 18842
rect 4140 18366 4158 18842
rect 4140 18362 4176 18366
rect 4072 18350 4176 18362
rect 3912 17580 3918 18060
rect 3974 17580 3982 18060
rect 3912 16328 3982 17580
rect 3912 15848 3924 16328
rect 3980 15848 3982 16328
rect 3912 14548 3982 15848
rect 3912 14068 3924 14548
rect 3980 14068 3982 14548
rect 3912 12914 3982 14068
rect 3912 12434 3914 12914
rect 3970 12434 3982 12914
rect 3912 11900 3982 12434
rect 4082 17208 4176 18350
rect 4082 16728 4090 17208
rect 4146 16728 4176 17208
rect 4082 15474 4176 16728
rect 4138 14994 4176 15474
rect 4082 13690 4176 14994
rect 4082 13210 4086 13690
rect 4142 13210 4176 13690
rect 4082 11902 4176 13210
rect 4530 18060 4600 19176
rect 4688 18852 4774 19896
rect 5140 19676 5210 19878
rect 5760 19676 5830 19878
rect 5136 19664 5220 19676
rect 5136 19184 5144 19664
rect 5136 19176 5220 19184
rect 5746 19664 5830 19676
rect 5746 19184 5754 19664
rect 5746 19176 5830 19184
rect 4688 18446 4702 18852
rect 4684 18372 4702 18446
rect 4758 18446 4774 18852
rect 4758 18372 4786 18446
rect 4684 18334 4786 18372
rect 4688 18330 4786 18334
rect 4530 17580 4538 18060
rect 4594 17580 4600 18060
rect 4530 16318 4600 17580
rect 4530 15838 4532 16318
rect 4588 15838 4600 16318
rect 4530 14550 4600 15838
rect 4530 14070 4532 14550
rect 4588 14070 4600 14550
rect 4530 12914 4600 14070
rect 4530 12434 4534 12914
rect 4590 12434 4600 12914
rect 4530 11902 4600 12434
rect 4692 17204 4786 18330
rect 4692 16724 4708 17204
rect 4764 16724 4786 17204
rect 4692 15486 4786 16724
rect 4692 15006 4704 15486
rect 4760 15006 4786 15486
rect 4692 13690 4786 15006
rect 4692 13210 4704 13690
rect 4760 13210 4786 13690
rect 4692 11902 4786 13210
rect 5140 18060 5210 19176
rect 5308 18848 5392 18918
rect 5308 18792 5320 18848
rect 5376 18792 5392 18848
rect 5140 17580 5148 18060
rect 5204 17580 5210 18060
rect 5140 16330 5210 17580
rect 5140 15850 5148 16330
rect 5204 15850 5210 16330
rect 5140 14542 5210 15850
rect 5140 14062 5148 14542
rect 5204 14062 5210 14542
rect 5140 12916 5210 14062
rect 5140 12436 5152 12916
rect 5208 12436 5210 12916
rect 5140 11902 5210 12436
rect 5302 18366 5382 18372
rect 5302 17210 5396 18366
rect 5302 16730 5310 17210
rect 5366 16730 5396 17210
rect 5302 15480 5396 16730
rect 5302 15000 5310 15480
rect 5366 15000 5396 15480
rect 5302 13694 5396 15000
rect 5358 13214 5396 13694
rect 5302 11902 5396 13214
rect 5760 18060 5830 19176
rect 5760 17580 5768 18060
rect 5824 17580 5830 18060
rect 5760 16320 5830 17580
rect 5760 15840 5774 16320
rect 5760 14544 5830 15840
rect 5760 14064 5766 14544
rect 5822 14064 5830 14544
rect 5760 12916 5830 14064
rect 5760 12436 5768 12916
rect 5824 12436 5830 12916
rect 5760 11902 5830 12436
rect 5912 18856 5990 19910
rect 6380 19674 6450 19878
rect 6348 19664 6450 19674
rect 6348 19184 6384 19664
rect 6440 19184 6450 19664
rect 6348 19174 6450 19184
rect 5912 18376 5932 18856
rect 5988 18376 5990 18856
rect 5912 18366 5990 18376
rect 5912 17206 6006 18366
rect 5912 16726 5920 17206
rect 5976 16726 6006 17206
rect 5912 15480 6006 16726
rect 5912 15000 5928 15480
rect 5984 15000 6006 15480
rect 5912 13692 6006 15000
rect 5912 13212 5926 13692
rect 5982 13212 6006 13692
rect 5912 11902 6006 13212
rect 6380 18060 6450 19174
rect 6516 18870 6594 19906
rect 6992 19676 7062 19872
rect 6992 19664 7078 19676
rect 6992 19184 7004 19664
rect 7060 19184 7078 19664
rect 6992 19176 7078 19184
rect 6516 18844 6620 18870
rect 6516 18368 6548 18844
rect 6604 18832 6620 18844
rect 6516 18366 6612 18368
rect 6516 18358 6616 18366
rect 6380 17580 6388 18060
rect 6444 17580 6450 18060
rect 6380 16330 6450 17580
rect 6380 15850 6386 16330
rect 6442 15850 6450 16330
rect 6380 14544 6450 15850
rect 6380 14064 6382 14544
rect 6438 14064 6450 14544
rect 6380 12928 6450 14064
rect 6380 12448 6390 12928
rect 6446 12448 6450 12928
rect 6380 11902 6450 12448
rect 6522 17202 6616 18358
rect 6522 16722 6540 17202
rect 6596 16722 6616 17202
rect 6522 15484 6616 16722
rect 6522 15004 6540 15484
rect 6596 15004 6616 15484
rect 6522 13696 6616 15004
rect 6522 13216 6540 13696
rect 6596 13216 6616 13696
rect 6522 11902 6616 13216
rect 6992 18060 7062 19176
rect 7140 18848 7236 19902
rect 7612 19678 7682 19872
rect 7608 19664 7692 19678
rect 7608 19184 7624 19664
rect 7680 19184 7692 19664
rect 7608 19178 7692 19184
rect 7140 18368 7166 18848
rect 7222 18368 7236 18848
rect 7140 18326 7236 18368
rect 6992 17580 6998 18060
rect 7054 17580 7062 18060
rect 6992 16324 7062 17580
rect 6992 15844 6996 16324
rect 7052 15844 7062 16324
rect 6992 14542 7062 15844
rect 6992 14062 7006 14542
rect 6992 12922 7062 14062
rect 6992 12442 7004 12922
rect 7060 12442 7062 12922
rect 6992 11896 7062 12442
rect 7142 17198 7236 18326
rect 7142 16718 7160 17198
rect 7216 16718 7236 17198
rect 7142 15488 7236 16718
rect 7142 15008 7158 15488
rect 7214 15008 7236 15488
rect 7142 13686 7236 15008
rect 7142 13206 7158 13686
rect 7214 13206 7236 13686
rect 7142 11902 7236 13206
rect 7612 18060 7682 19178
rect 7612 17580 7618 18060
rect 7674 17580 7682 18060
rect 7612 16326 7682 17580
rect 7612 15846 7624 16326
rect 7680 15846 7682 16326
rect 7612 14544 7682 15846
rect 7612 14064 7624 14544
rect 7680 14064 7682 14544
rect 7612 12922 7682 14064
rect 7612 12442 7622 12922
rect 7678 12442 7682 12922
rect 7612 11896 7682 12442
rect 7752 18850 7862 19906
rect 8232 19680 8302 19872
rect 8230 19664 8314 19680
rect 8230 19184 8244 19664
rect 8300 19184 8314 19664
rect 8230 19180 8314 19184
rect 7752 18370 7780 18850
rect 7836 18370 7862 18850
rect 7752 18326 7862 18370
rect 7752 17194 7846 18326
rect 7752 16714 7774 17194
rect 7830 16714 7846 17194
rect 7752 15474 7846 16714
rect 7752 14994 7760 15474
rect 7816 14994 7846 15474
rect 7752 13696 7846 14994
rect 7752 13216 7776 13696
rect 7832 13216 7846 13696
rect 7752 11902 7846 13216
rect 8232 18060 8302 19180
rect 8366 18850 8476 19900
rect 8842 19678 8912 19872
rect 8836 19664 8920 19678
rect 9452 19674 9522 19872
rect 10072 19674 10142 19872
rect 10692 19676 10762 19872
rect 8836 19184 8854 19664
rect 8910 19184 8920 19664
rect 8836 19178 8920 19184
rect 9446 19664 9530 19674
rect 9446 19184 9464 19664
rect 9520 19184 9530 19664
rect 8366 18400 8396 18850
rect 8356 18370 8396 18400
rect 8452 18370 8476 18850
rect 8356 18354 8476 18370
rect 8232 17580 8238 18060
rect 8294 17580 8302 18060
rect 8232 16326 8302 17580
rect 8232 15846 8240 16326
rect 8296 15846 8302 16326
rect 8232 14544 8302 15846
rect 8232 14064 8236 14544
rect 8292 14064 8302 14544
rect 8232 12920 8302 14064
rect 8288 12440 8302 12920
rect 8232 11896 8302 12440
rect 8362 18320 8476 18354
rect 8362 17198 8456 18320
rect 8362 16718 8390 17198
rect 8446 16718 8456 17198
rect 8362 15476 8456 16718
rect 8362 14996 8390 15476
rect 8446 14996 8456 15476
rect 8362 13700 8456 14996
rect 8362 13220 8394 13700
rect 8450 13220 8456 13700
rect 8362 11902 8456 13220
rect 8842 18060 8912 19178
rect 9446 19174 9530 19184
rect 10070 19664 10154 19674
rect 10070 19184 10084 19664
rect 10140 19184 10154 19664
rect 10070 19174 10154 19184
rect 10688 19664 10772 19676
rect 11312 19674 11382 19872
rect 11932 19676 12002 19872
rect 12542 19678 12612 19872
rect 10688 19184 10704 19664
rect 10760 19184 10772 19664
rect 10688 19176 10772 19184
rect 11300 19664 11384 19674
rect 11300 19184 11314 19664
rect 11370 19184 11384 19664
rect 8842 17580 8848 18060
rect 8904 17580 8912 18060
rect 8842 16320 8912 17580
rect 8842 15840 8852 16320
rect 8908 15840 8912 16320
rect 8842 14542 8912 15840
rect 8842 14062 8856 14542
rect 8842 12918 8912 14062
rect 8842 12438 8854 12918
rect 8910 12438 8912 12918
rect 8842 11896 8912 12438
rect 8982 18850 9094 18894
rect 8982 18370 9016 18850
rect 9072 18370 9094 18850
rect 8982 18318 9094 18370
rect 8982 17202 9076 18318
rect 8982 16722 9010 17202
rect 9066 16722 9076 17202
rect 8982 15484 9076 16722
rect 8982 15004 9004 15484
rect 9060 15004 9076 15484
rect 8982 13700 9076 15004
rect 8982 13220 9000 13700
rect 9056 13220 9076 13700
rect 8982 11902 9076 13220
rect 9452 18060 9522 19174
rect 9608 18850 9724 18862
rect 9608 18370 9624 18850
rect 9680 18370 9724 18850
rect 9608 18324 9724 18370
rect 9452 17580 9458 18060
rect 9514 17580 9522 18060
rect 9452 16316 9522 17580
rect 9452 15836 9466 16316
rect 9452 14542 9522 15836
rect 9452 14062 9466 14542
rect 9452 12916 9522 14062
rect 9452 12436 9466 12916
rect 9452 11896 9522 12436
rect 9612 17202 9706 18324
rect 9612 16722 9624 17202
rect 9680 16722 9706 17202
rect 9612 15476 9706 16722
rect 9612 14996 9632 15476
rect 9688 14996 9706 15476
rect 9612 13692 9706 14996
rect 9612 13212 9622 13692
rect 9678 13212 9706 13692
rect 9612 11902 9706 13212
rect 10072 18060 10142 19174
rect 10236 18854 10352 18866
rect 10236 18374 10246 18854
rect 10302 18374 10352 18854
rect 10236 18328 10352 18374
rect 10072 17580 10078 18060
rect 10134 17580 10142 18060
rect 10072 16326 10142 17580
rect 10072 15846 10078 16326
rect 10134 15846 10142 16326
rect 10242 17198 10336 18328
rect 10242 16718 10246 17198
rect 10302 16718 10336 17198
rect 10242 16322 10336 16718
rect 10072 14536 10142 15846
rect 10236 15840 10336 16322
rect 10072 14056 10076 14536
rect 10132 14056 10142 14536
rect 10072 12926 10142 14056
rect 10072 12446 10082 12926
rect 10138 12446 10142 12926
rect 10072 11896 10142 12446
rect 10242 15478 10336 15840
rect 10242 14998 10248 15478
rect 10304 14998 10336 15478
rect 10242 13692 10336 14998
rect 10242 13212 10244 13692
rect 10300 13212 10336 13692
rect 10242 11902 10336 13212
rect 10692 18060 10762 19176
rect 11300 19174 11384 19184
rect 11916 19664 12002 19676
rect 11916 19184 11934 19664
rect 11990 19184 12002 19664
rect 11916 19176 12002 19184
rect 12534 19664 12618 19678
rect 13152 19676 13222 19872
rect 13772 19676 13842 19872
rect 12534 19184 12554 19664
rect 12610 19184 12618 19664
rect 12534 19178 12618 19184
rect 13150 19664 13234 19676
rect 13150 19184 13164 19664
rect 13220 19184 13234 19664
rect 10848 18848 10976 18858
rect 10848 18368 10856 18848
rect 10912 18368 10976 18848
rect 10848 18330 10976 18368
rect 10692 17580 10698 18060
rect 10754 17580 10762 18060
rect 10692 16328 10762 17580
rect 10692 15848 10702 16328
rect 10758 15848 10762 16328
rect 10692 14540 10762 15848
rect 10692 14060 10704 14540
rect 10760 14060 10762 14540
rect 10692 12918 10762 14060
rect 10692 12438 10694 12918
rect 10750 12438 10762 12918
rect 10692 11896 10762 12438
rect 10862 17200 10956 18330
rect 10918 16720 10956 17200
rect 10862 15486 10956 16720
rect 10918 15006 10956 15486
rect 10862 13690 10956 15006
rect 10862 13210 10866 13690
rect 10922 13210 10956 13690
rect 10862 11902 10956 13210
rect 11312 18060 11382 19174
rect 11464 18850 11592 18860
rect 11464 18370 11476 18850
rect 11532 18370 11592 18850
rect 11464 18332 11592 18370
rect 11312 17580 11318 18060
rect 11374 17580 11382 18060
rect 11312 16324 11382 17580
rect 11312 15844 11320 16324
rect 11376 15844 11382 16324
rect 11312 14540 11382 15844
rect 11312 14060 11314 14540
rect 11370 14060 11382 14540
rect 11312 12916 11382 14060
rect 11312 12436 11316 12916
rect 11372 12436 11382 12916
rect 11312 11896 11382 12436
rect 11472 17198 11566 18332
rect 11472 16718 11476 17198
rect 11532 16718 11566 17198
rect 11472 15482 11566 16718
rect 11472 15002 11480 15482
rect 11536 15002 11566 15482
rect 11472 13692 11566 15002
rect 11472 13212 11484 13692
rect 11540 13212 11566 13692
rect 11472 11902 11566 13212
rect 11932 18060 12002 19176
rect 12064 18848 12192 18856
rect 12064 18368 12092 18848
rect 12148 18368 12192 18848
rect 12064 18328 12192 18368
rect 11932 17580 11938 18060
rect 11994 17580 12002 18060
rect 11932 16324 12002 17580
rect 11932 15844 11940 16324
rect 11996 15844 12002 16324
rect 11932 14544 12002 15844
rect 11932 14064 11940 14544
rect 11996 14064 12002 14544
rect 11932 12918 12002 14064
rect 11932 12438 11938 12918
rect 11994 12438 12002 12918
rect 11932 11896 12002 12438
rect 12082 17210 12176 18328
rect 12082 16730 12096 17210
rect 12152 16730 12176 17210
rect 12082 15486 12176 16730
rect 12082 15006 12094 15486
rect 12150 15006 12176 15486
rect 12082 13692 12176 15006
rect 12082 13212 12094 13692
rect 12150 13212 12176 13692
rect 12082 11902 12176 13212
rect 12542 18060 12612 19178
rect 13150 19176 13234 19184
rect 13750 19664 13842 19676
rect 13750 19184 13774 19664
rect 13830 19184 13842 19664
rect 13750 19176 13842 19184
rect 12692 18850 12820 18864
rect 12692 18370 12712 18850
rect 12768 18370 12820 18850
rect 12692 18336 12820 18370
rect 12542 17580 12548 18060
rect 12604 17580 12612 18060
rect 12542 16316 12612 17580
rect 12542 15836 12550 16316
rect 12606 15836 12612 16316
rect 12542 14540 12612 15836
rect 12542 14060 12554 14540
rect 12610 14060 12612 14540
rect 12542 12926 12612 14060
rect 12542 12446 12550 12926
rect 12606 12446 12612 12926
rect 12542 11896 12612 12446
rect 12702 17198 12796 18336
rect 12758 16718 12796 17198
rect 12702 15482 12796 16718
rect 12702 15002 12718 15482
rect 12774 15002 12796 15482
rect 12702 13686 12796 15002
rect 12702 13206 12710 13686
rect 12766 13206 12796 13686
rect 12702 11902 12796 13206
rect 13152 18060 13222 19176
rect 13298 18856 13426 18868
rect 13298 18376 13322 18856
rect 13378 18376 13426 18856
rect 13298 18340 13426 18376
rect 13152 17580 13158 18060
rect 13214 17580 13222 18060
rect 13152 16320 13222 17580
rect 13152 15840 13162 16320
rect 13218 15840 13222 16320
rect 13152 14540 13222 15840
rect 13152 14060 13162 14540
rect 13218 14060 13222 14540
rect 13152 12924 13222 14060
rect 13152 12444 13164 12924
rect 13220 12444 13222 12924
rect 13152 11896 13222 12444
rect 13312 17206 13406 18340
rect 13312 16726 13316 17206
rect 13372 16726 13406 17206
rect 13312 15486 13406 16726
rect 13312 15006 13314 15486
rect 13370 15006 13406 15486
rect 13312 13688 13406 15006
rect 13312 13208 13324 13688
rect 13380 13208 13406 13688
rect 13312 11902 13406 13208
rect 13772 18060 13842 19176
rect 13904 18844 14032 18858
rect 13904 18368 13940 18844
rect 13996 18368 14032 18844
rect 13904 18330 14032 18368
rect 13772 17580 13778 18060
rect 13834 17580 13842 18060
rect 13772 16324 13842 17580
rect 13772 15844 13778 16324
rect 13834 15844 13842 16324
rect 13772 14538 13842 15844
rect 13772 14058 13786 14538
rect 13772 12922 13842 14058
rect 13772 12442 13784 12922
rect 13840 12442 13842 12922
rect 13772 11896 13842 12442
rect 13922 17198 14016 18330
rect 13922 16718 13940 17198
rect 13996 16718 14016 17198
rect 13922 15486 14016 16718
rect 13922 15006 13932 15486
rect 13988 15006 14016 15486
rect 13922 13694 14016 15006
rect 13922 13214 13940 13694
rect 13996 13214 14016 13694
rect 13922 11902 14016 13214
rect 2118 11750 14048 11860
<< via1 >>
rect 2084 19184 2140 19664
rect 2072 17568 2128 18048
rect 2066 15846 2122 16326
rect 2076 14064 2132 14544
rect 2066 12448 2122 12928
rect 2234 18366 2290 18846
rect 2236 16728 2292 17208
rect 2234 15008 2290 15488
rect 2226 13212 2282 13692
rect 2694 19184 2750 19664
rect 3304 19184 3360 19664
rect 2852 18364 2908 18844
rect 2688 17580 2744 18060
rect 2688 15842 2744 16322
rect 2688 14068 2744 14548
rect 2688 12438 2744 12918
rect 2852 16714 2908 17194
rect 2854 14994 2910 15474
rect 2848 13206 2904 13686
rect 3924 19184 3980 19664
rect 3470 18372 3526 18852
rect 3308 17580 3364 18060
rect 3312 15846 3368 16326
rect 3308 14064 3364 14544
rect 3308 12446 3364 12926
rect 3478 16730 3534 17210
rect 3474 15008 3530 15488
rect 3470 13220 3526 13700
rect 4534 19184 4600 19664
rect 4084 18362 4140 18842
rect 3918 17580 3974 18060
rect 3924 15848 3980 16328
rect 3924 14068 3980 14548
rect 3914 12434 3970 12914
rect 4090 16728 4146 17208
rect 4082 14994 4138 15474
rect 4086 13210 4142 13690
rect 5144 19184 5220 19664
rect 5754 19184 5830 19664
rect 4702 18372 4758 18852
rect 4538 17580 4594 18060
rect 4532 15838 4588 16318
rect 4532 14070 4588 14550
rect 4534 12434 4590 12914
rect 4708 16724 4764 17204
rect 4704 15006 4760 15486
rect 4704 13210 4760 13690
rect 5320 18372 5376 18848
rect 5148 17580 5204 18060
rect 5148 15850 5204 16330
rect 5148 14062 5204 14542
rect 5152 12436 5208 12916
rect 5310 16730 5366 17210
rect 5310 15000 5366 15480
rect 5302 13214 5358 13694
rect 5768 17580 5824 18060
rect 5774 15840 5830 16320
rect 5766 14064 5822 14544
rect 5768 12436 5824 12916
rect 6384 19184 6440 19664
rect 5932 18376 5988 18856
rect 5920 16726 5976 17206
rect 5928 15000 5984 15480
rect 5926 13212 5982 13692
rect 7004 19184 7060 19664
rect 6548 18368 6604 18844
rect 6388 17580 6444 18060
rect 6386 15850 6442 16330
rect 6382 14064 6438 14544
rect 6390 12448 6446 12928
rect 6540 16722 6596 17202
rect 6540 15004 6596 15484
rect 6540 13216 6596 13696
rect 7624 19184 7680 19664
rect 7166 18368 7222 18848
rect 6998 17580 7054 18060
rect 6996 15844 7052 16324
rect 7006 14062 7062 14542
rect 7004 12442 7060 12922
rect 7160 16718 7216 17198
rect 7158 15008 7214 15488
rect 7158 13206 7214 13686
rect 7618 17580 7674 18060
rect 7624 15846 7680 16326
rect 7624 14064 7680 14544
rect 7622 12442 7678 12922
rect 8244 19184 8300 19664
rect 7780 18370 7836 18850
rect 7774 16714 7830 17194
rect 7760 14994 7816 15474
rect 7776 13216 7832 13696
rect 8854 19184 8910 19664
rect 9464 19184 9520 19664
rect 8396 18370 8452 18850
rect 8238 17580 8294 18060
rect 8240 15846 8296 16326
rect 8236 14064 8292 14544
rect 8232 12440 8288 12920
rect 8390 16718 8446 17198
rect 8390 14996 8446 15476
rect 8394 13220 8450 13700
rect 10084 19184 10140 19664
rect 10704 19184 10760 19664
rect 11314 19184 11370 19664
rect 8848 17580 8904 18060
rect 8852 15840 8908 16320
rect 8856 14062 8912 14542
rect 8854 12438 8910 12918
rect 9016 18370 9072 18850
rect 9010 16722 9066 17202
rect 9004 15004 9060 15484
rect 9000 13220 9056 13700
rect 9624 18370 9680 18850
rect 9458 17580 9514 18060
rect 9466 15836 9522 16316
rect 9466 14062 9522 14542
rect 9466 12436 9522 12916
rect 9624 16722 9680 17202
rect 9632 14996 9688 15476
rect 9622 13212 9678 13692
rect 10246 18374 10302 18854
rect 10078 17580 10134 18060
rect 10078 15846 10134 16326
rect 10246 16718 10302 17198
rect 10076 14056 10132 14536
rect 10082 12446 10138 12926
rect 10248 14998 10304 15478
rect 10244 13212 10300 13692
rect 11934 19184 11990 19664
rect 12554 19184 12610 19664
rect 13164 19184 13220 19664
rect 10856 18368 10912 18848
rect 10698 17580 10754 18060
rect 10702 15848 10758 16328
rect 10704 14060 10760 14540
rect 10694 12438 10750 12918
rect 10862 16720 10918 17200
rect 10862 15006 10918 15486
rect 10866 13210 10922 13690
rect 11476 18370 11532 18850
rect 11318 17580 11374 18060
rect 11320 15844 11376 16324
rect 11314 14060 11370 14540
rect 11316 12436 11372 12916
rect 11476 16718 11532 17198
rect 11480 15002 11536 15482
rect 11484 13212 11540 13692
rect 12092 18368 12148 18848
rect 11938 17580 11994 18060
rect 11940 15844 11996 16324
rect 11940 14064 11996 14544
rect 11938 12438 11994 12918
rect 12096 16730 12152 17210
rect 12094 15006 12150 15486
rect 12094 13212 12150 13692
rect 13774 19184 13830 19664
rect 12712 18370 12768 18850
rect 12548 17580 12604 18060
rect 12550 15836 12606 16316
rect 12554 14060 12610 14540
rect 12550 12446 12606 12926
rect 12702 16718 12758 17198
rect 12718 15002 12774 15482
rect 12710 13206 12766 13686
rect 13322 18376 13378 18856
rect 13158 17580 13214 18060
rect 13162 15840 13218 16320
rect 13162 14060 13218 14540
rect 13164 12444 13220 12924
rect 13316 16726 13372 17206
rect 13314 15006 13370 15486
rect 13324 13208 13380 13688
rect 13940 18368 13996 18844
rect 13778 17580 13834 18060
rect 13778 15844 13834 16324
rect 13786 14058 13842 14538
rect 13784 12442 13840 12922
rect 13940 16718 13996 17198
rect 13932 15006 13988 15486
rect 13940 13214 13996 13694
<< metal2 >>
rect 14378 20706 14806 20746
rect 13676 20642 14806 20706
rect 1242 19676 1662 20194
rect 14378 20112 14806 20642
rect 1242 19674 1892 19676
rect 6516 19674 6594 19906
rect 14378 19872 14804 20112
rect 1242 19664 14204 19674
rect 1242 19184 2084 19664
rect 2140 19184 2694 19664
rect 2750 19184 3304 19664
rect 3360 19184 3924 19664
rect 3980 19184 4534 19664
rect 4600 19184 5144 19664
rect 5220 19184 5754 19664
rect 5830 19184 6384 19664
rect 6440 19184 7004 19664
rect 7060 19184 7624 19664
rect 7680 19184 8244 19664
rect 8300 19184 8854 19664
rect 8910 19184 9464 19664
rect 9520 19184 10084 19664
rect 10140 19184 10704 19664
rect 10760 19184 11314 19664
rect 11370 19184 11934 19664
rect 11990 19184 12554 19664
rect 12610 19184 13164 19664
rect 13220 19184 13774 19664
rect 13830 19184 14204 19664
rect 1242 19178 14204 19184
rect 1242 19176 1892 19178
rect 1242 18064 1662 19176
rect 14380 18858 14800 19872
rect 14198 18856 14800 18858
rect 1874 18852 5932 18856
rect 1874 18846 3470 18852
rect 1874 18366 2234 18846
rect 2290 18844 3470 18846
rect 2290 18366 2852 18844
rect 1874 18364 2852 18366
rect 2908 18372 3470 18844
rect 3526 18842 4702 18852
rect 3526 18372 4084 18842
rect 2908 18364 4084 18372
rect 1874 18362 4084 18364
rect 4140 18372 4702 18842
rect 4758 18848 5932 18852
rect 4758 18372 5320 18848
rect 5376 18376 5932 18848
rect 5988 18854 13322 18856
rect 5988 18850 10246 18854
rect 5988 18848 7780 18850
rect 5988 18844 7166 18848
rect 5988 18376 6548 18844
rect 5376 18372 6548 18376
rect 4140 18368 6548 18372
rect 6604 18368 7166 18844
rect 7222 18370 7780 18848
rect 7836 18370 8396 18850
rect 8452 18370 9016 18850
rect 9072 18370 9624 18850
rect 9680 18374 10246 18850
rect 10302 18850 13322 18854
rect 10302 18848 11476 18850
rect 10302 18374 10856 18848
rect 9680 18370 10856 18374
rect 7222 18368 10856 18370
rect 10912 18370 11476 18848
rect 11532 18848 12712 18850
rect 11532 18370 12092 18848
rect 10912 18368 12092 18370
rect 12148 18370 12712 18848
rect 12768 18376 13322 18850
rect 13378 18844 14800 18856
rect 13378 18376 13940 18844
rect 12768 18370 13940 18376
rect 12148 18368 13940 18370
rect 13996 18368 14800 18844
rect 4140 18364 14800 18368
rect 4140 18362 5912 18364
rect 1874 18360 5912 18362
rect 5980 18360 14800 18364
rect 4684 18334 4786 18360
rect 6516 18358 6594 18360
rect 14198 18358 14800 18360
rect 1242 18062 1920 18064
rect 1242 18060 14202 18062
rect 1242 18048 2688 18060
rect 1242 17568 2072 18048
rect 2128 17580 2688 18048
rect 2744 17580 3308 18060
rect 3364 17580 3918 18060
rect 3974 17580 4538 18060
rect 4594 17580 5148 18060
rect 5204 17580 5768 18060
rect 5824 17580 6388 18060
rect 6444 17580 6998 18060
rect 7054 17580 7618 18060
rect 7674 17580 8238 18060
rect 8294 17580 8848 18060
rect 8904 17580 9458 18060
rect 9514 17580 10078 18060
rect 10134 17580 10698 18060
rect 10754 17580 11318 18060
rect 11374 17580 11938 18060
rect 11994 17580 12548 18060
rect 12604 17580 13158 18060
rect 13214 17580 13778 18060
rect 13834 17580 14202 18060
rect 2128 17568 14202 17580
rect 1242 17566 14202 17568
rect 1242 17564 1920 17566
rect 1242 16332 1662 17564
rect 14380 17214 14800 18358
rect 14202 17210 14800 17214
rect 1874 17208 3478 17210
rect 1874 16728 2236 17208
rect 2292 17194 3478 17208
rect 2292 16728 2852 17194
rect 1874 16714 2852 16728
rect 2908 16730 3478 17194
rect 3534 17208 5310 17210
rect 3534 16730 4090 17208
rect 2908 16728 4090 16730
rect 4146 17204 5310 17208
rect 4146 16728 4708 17204
rect 2908 16724 4708 16728
rect 4764 16730 5310 17204
rect 5366 17206 12096 17210
rect 5366 16730 5920 17206
rect 4764 16726 5920 16730
rect 5976 17202 12096 17206
rect 5976 16726 6540 17202
rect 4764 16724 6540 16726
rect 2908 16722 6540 16724
rect 6596 17198 9010 17202
rect 6596 16722 7160 17198
rect 2908 16718 7160 16722
rect 7216 17194 8390 17198
rect 7216 16718 7774 17194
rect 2908 16714 7774 16718
rect 7830 16718 8390 17194
rect 8446 16722 9010 17198
rect 9066 16722 9624 17202
rect 9680 17200 12096 17202
rect 9680 17198 10862 17200
rect 9680 16722 10246 17198
rect 8446 16718 10246 16722
rect 10302 16720 10862 17198
rect 10918 17198 12096 17200
rect 10918 16720 11476 17198
rect 10302 16718 11476 16720
rect 11532 16730 12096 17198
rect 12152 17206 14800 17210
rect 12152 17198 13316 17206
rect 12152 16730 12702 17198
rect 11532 16718 12702 16730
rect 12758 16726 13316 17198
rect 13372 17198 14800 17206
rect 13372 16726 13940 17198
rect 12758 16718 13940 16726
rect 13996 16718 14800 17198
rect 7830 16714 14800 16718
rect 1242 16330 1922 16332
rect 1242 16328 5148 16330
rect 1242 16326 3924 16328
rect 1242 15846 2066 16326
rect 2122 16322 3312 16326
rect 2122 15846 2688 16322
rect 1242 15842 2688 15846
rect 2744 15846 3312 16322
rect 3368 15848 3924 16326
rect 3980 16318 5148 16328
rect 3980 15848 4532 16318
rect 3368 15846 4532 15848
rect 2744 15842 4532 15846
rect 1242 15838 4532 15842
rect 4588 15850 5148 16318
rect 5204 16320 6386 16330
rect 5204 15850 5774 16320
rect 4588 15840 5774 15850
rect 5830 15850 6386 16320
rect 6442 16328 14212 16330
rect 6442 16326 10702 16328
rect 6442 16324 7624 16326
rect 6442 15850 6996 16324
rect 5830 15844 6996 15850
rect 7052 15846 7624 16324
rect 7680 15846 8240 16326
rect 8296 16320 10078 16326
rect 8296 15846 8852 16320
rect 7052 15844 8852 15846
rect 5830 15840 8852 15844
rect 8908 16316 10078 16320
rect 8908 15840 9466 16316
rect 4588 15838 9466 15840
rect 1242 15836 9466 15838
rect 9522 15846 10078 16316
rect 10134 15848 10702 16326
rect 10758 16324 14212 16328
rect 10758 15848 11320 16324
rect 10134 15846 11320 15848
rect 9522 15844 11320 15846
rect 11376 15844 11940 16324
rect 11996 16320 13778 16324
rect 11996 16316 13162 16320
rect 11996 15844 12550 16316
rect 9522 15836 12550 15844
rect 12606 15840 13162 16316
rect 13218 15844 13778 16320
rect 13834 15844 14212 16324
rect 13218 15840 14212 15844
rect 12606 15836 14212 15840
rect 1242 15834 14212 15836
rect 1242 15832 1922 15834
rect 1242 14550 1662 15832
rect 14380 15488 14800 16714
rect 1876 15008 2234 15488
rect 2290 15474 3474 15488
rect 2290 15008 2854 15474
rect 1876 14994 2854 15008
rect 2910 15008 3474 15474
rect 3530 15486 7158 15488
rect 3530 15474 4704 15486
rect 3530 15008 4082 15474
rect 2910 14994 4082 15008
rect 4138 15006 4704 15474
rect 4760 15484 7158 15486
rect 4760 15480 6540 15484
rect 4760 15006 5310 15480
rect 4138 15000 5310 15006
rect 5366 15000 5928 15480
rect 5984 15004 6540 15480
rect 6596 15008 7158 15484
rect 7214 15486 14800 15488
rect 7214 15484 10862 15486
rect 7214 15476 9004 15484
rect 7214 15474 8390 15476
rect 7214 15008 7760 15474
rect 6596 15004 7760 15008
rect 5984 15000 7760 15004
rect 4138 14994 7760 15000
rect 7816 14996 8390 15474
rect 8446 15004 9004 15476
rect 9060 15478 10862 15484
rect 9060 15476 10248 15478
rect 9060 15004 9632 15476
rect 8446 14996 9632 15004
rect 9688 14998 10248 15476
rect 10304 15006 10862 15478
rect 10918 15482 12094 15486
rect 10918 15006 11480 15482
rect 10304 15002 11480 15006
rect 11536 15006 12094 15482
rect 12150 15482 13314 15486
rect 12150 15006 12718 15482
rect 11536 15002 12718 15006
rect 12774 15006 13314 15482
rect 13370 15006 13932 15486
rect 13988 15006 14800 15486
rect 12774 15002 14800 15006
rect 10304 14998 14800 15002
rect 9688 14996 14800 14998
rect 7816 14994 14800 14996
rect 1876 14992 14800 14994
rect 14206 14988 14800 14992
rect 1242 14548 4532 14550
rect 1242 14544 2688 14548
rect 1242 14064 2076 14544
rect 2132 14068 2688 14544
rect 2744 14544 3924 14548
rect 2744 14068 3308 14544
rect 2132 14064 3308 14068
rect 3364 14068 3924 14544
rect 3980 14070 4532 14548
rect 4588 14544 14200 14550
rect 4588 14542 5766 14544
rect 4588 14070 5148 14542
rect 3980 14068 5148 14070
rect 3364 14064 5148 14068
rect 1242 14062 5148 14064
rect 5204 14064 5766 14542
rect 5822 14064 6382 14544
rect 6438 14542 7624 14544
rect 6438 14064 7006 14542
rect 5204 14062 7006 14064
rect 7062 14064 7624 14542
rect 7680 14064 8236 14544
rect 8292 14542 11940 14544
rect 8292 14064 8856 14542
rect 7062 14062 8856 14064
rect 8912 14062 9466 14542
rect 9522 14540 11940 14542
rect 9522 14536 10704 14540
rect 9522 14062 10076 14536
rect 1242 14056 10076 14062
rect 10132 14060 10704 14536
rect 10760 14060 11314 14540
rect 11370 14064 11940 14540
rect 11996 14540 14200 14544
rect 11996 14064 12554 14540
rect 11370 14060 12554 14064
rect 12610 14060 13162 14540
rect 13218 14538 14200 14540
rect 13218 14060 13786 14538
rect 10132 14058 13786 14060
rect 13842 14058 14200 14538
rect 10132 14056 14200 14058
rect 1242 13724 1662 14056
rect 1864 14054 14200 14056
rect 1242 13198 1660 13724
rect 14380 13704 14800 14988
rect 14206 13700 14800 13704
rect 1878 13692 3470 13700
rect 1878 13212 2226 13692
rect 2282 13686 3470 13692
rect 2282 13212 2848 13686
rect 1878 13206 2848 13212
rect 2904 13220 3470 13686
rect 3526 13696 8394 13700
rect 3526 13694 6540 13696
rect 3526 13690 5302 13694
rect 3526 13220 4086 13690
rect 2904 13210 4086 13220
rect 4142 13210 4704 13690
rect 4760 13214 5302 13690
rect 5358 13692 6540 13694
rect 5358 13214 5926 13692
rect 4760 13212 5926 13214
rect 5982 13216 6540 13692
rect 6596 13686 7776 13696
rect 6596 13216 7158 13686
rect 5982 13212 7158 13216
rect 4760 13210 7158 13212
rect 2904 13206 7158 13210
rect 7214 13216 7776 13686
rect 7832 13220 8394 13696
rect 8450 13220 9000 13700
rect 9056 13694 14800 13700
rect 9056 13692 13940 13694
rect 9056 13220 9622 13692
rect 7832 13216 9622 13220
rect 7214 13212 9622 13216
rect 9678 13212 10244 13692
rect 10300 13690 11484 13692
rect 10300 13212 10866 13690
rect 7214 13210 10866 13212
rect 10922 13212 11484 13690
rect 11540 13212 12094 13692
rect 12150 13688 13940 13692
rect 12150 13686 13324 13688
rect 12150 13212 12710 13686
rect 10922 13210 12710 13212
rect 7214 13206 12710 13210
rect 12766 13208 13324 13686
rect 13380 13214 13940 13688
rect 13996 13214 14800 13694
rect 13380 13208 14800 13214
rect 12766 13206 14800 13208
rect 1878 13204 14800 13206
rect 1242 12928 1662 13198
rect 1242 12448 2066 12928
rect 2122 12926 6390 12928
rect 2122 12918 3308 12926
rect 2122 12448 2688 12918
rect 1242 12438 2688 12448
rect 2744 12446 3308 12918
rect 3364 12916 6390 12926
rect 3364 12914 5152 12916
rect 3364 12446 3914 12914
rect 2744 12438 3914 12446
rect 1242 12434 3914 12438
rect 3970 12434 4534 12914
rect 4590 12436 5152 12914
rect 5208 12436 5768 12916
rect 5824 12448 6390 12916
rect 6446 12926 14208 12928
rect 6446 12922 10082 12926
rect 6446 12448 7004 12922
rect 5824 12442 7004 12448
rect 7060 12442 7622 12922
rect 7678 12920 10082 12922
rect 7678 12442 8232 12920
rect 5824 12440 8232 12442
rect 8288 12918 10082 12920
rect 8288 12440 8854 12918
rect 5824 12438 8854 12440
rect 8910 12916 10082 12918
rect 8910 12438 9466 12916
rect 5824 12436 9466 12438
rect 9522 12446 10082 12916
rect 10138 12918 12550 12926
rect 10138 12446 10694 12918
rect 9522 12438 10694 12446
rect 10750 12916 11938 12918
rect 10750 12438 11316 12916
rect 9522 12436 11316 12438
rect 11372 12438 11938 12916
rect 11994 12446 12550 12918
rect 12606 12924 14208 12926
rect 12606 12446 13164 12924
rect 11994 12444 13164 12446
rect 13220 12922 14208 12924
rect 13220 12444 13784 12922
rect 11994 12442 13784 12444
rect 13840 12442 14208 12922
rect 11994 12438 14208 12442
rect 11372 12436 14208 12438
rect 4590 12434 14208 12436
rect 1242 12432 14208 12434
rect 1242 11596 1662 12432
rect 14380 11610 14800 13204
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_0
timestamp 1666636516
transform 1 0 2185 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_1
timestamp 1666636516
transform 1 0 2801 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_2
timestamp 1666636516
transform 1 0 3417 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_3
timestamp 1666636516
transform 1 0 4033 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_4
timestamp 1666636516
transform 1 0 4649 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_5
timestamp 1666636516
transform 1 0 5265 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_6
timestamp 1666636516
transform 1 0 5881 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_7
timestamp 1666636516
transform 1 0 6497 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_8
timestamp 1666636516
transform 1 0 7113 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_9
timestamp 1666636516
transform 1 0 7729 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_10
timestamp 1666636516
transform 1 0 8345 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_11
timestamp 1666636516
transform 1 0 8961 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_12
timestamp 1666636516
transform 1 0 9577 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_13
timestamp 1666636516
transform 1 0 10193 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_14
timestamp 1666636516
transform 1 0 10809 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_15
timestamp 1666636516
transform 1 0 11425 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_16
timestamp 1666636516
transform 1 0 12041 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_17
timestamp 1666636516
transform 1 0 12657 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_18
timestamp 1666636516
transform 1 0 13273 0 1 15900
box -308 -4297 308 4297
use sky130_fd_pr__pfet_g5v0d10v5_WEH7DU  sky130_fd_pr__pfet_g5v0d10v5_WEH7DU_19
timestamp 1666636516
transform 1 0 13889 0 1 15900
box -308 -4297 308 4297
<< end >>
