magic
tech sky130A
timestamp 1665661005
<< metal4 >>
rect -675 -550 424 550
<< mimcap2 >>
rect -625 480 374 500
rect -625 -480 -605 480
rect 354 -480 374 480
rect -625 -500 374 -480
<< mimcap2contact >>
rect -605 -480 354 480
<< metal5 >>
rect -617 480 366 492
rect -617 -480 -605 480
rect 354 -480 366 480
rect -617 -492 366 -480
<< properties >>
string FIXED_BBOX -675 -550 424 550
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 10 l 10 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
