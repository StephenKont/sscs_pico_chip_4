magic
tech sky130A
magscale 1 2
timestamp 1668275587
<< pwell >>
rect -18850 29784 -3976 29936
rect -18850 13216 -18698 29784
rect -4128 13216 -3976 29784
rect -18850 13064 -3976 13216
<< psubdiff >>
rect -4060 29910 -4014 29916
rect -18824 29877 -4014 29910
rect -18824 29843 -18708 29877
rect -18674 29843 -18618 29877
rect -18584 29843 -18528 29877
rect -18494 29843 -18438 29877
rect -18404 29843 -18348 29877
rect -18314 29843 -18258 29877
rect -18224 29843 -18168 29877
rect -18134 29843 -18078 29877
rect -18044 29843 -17988 29877
rect -17954 29843 -17898 29877
rect -17864 29843 -17808 29877
rect -17774 29843 -17718 29877
rect -17684 29843 -17628 29877
rect -17594 29843 -17420 29877
rect -17386 29843 -17330 29877
rect -17296 29843 -17240 29877
rect -17206 29843 -17150 29877
rect -17116 29843 -17060 29877
rect -17026 29843 -16970 29877
rect -16936 29843 -16880 29877
rect -16846 29843 -16790 29877
rect -16756 29843 -16700 29877
rect -16666 29843 -16610 29877
rect -16576 29843 -16520 29877
rect -16486 29843 -16430 29877
rect -16396 29843 -16340 29877
rect -16306 29843 -16132 29877
rect -16098 29843 -16042 29877
rect -16008 29843 -15952 29877
rect -15918 29843 -15862 29877
rect -15828 29843 -15772 29877
rect -15738 29843 -15682 29877
rect -15648 29843 -15592 29877
rect -15558 29843 -15502 29877
rect -15468 29843 -15412 29877
rect -15378 29843 -15322 29877
rect -15288 29843 -15232 29877
rect -15198 29843 -15142 29877
rect -15108 29843 -15052 29877
rect -15018 29843 -14916 29877
rect -14882 29843 -14826 29877
rect -14792 29843 -14736 29877
rect -14702 29843 -14646 29877
rect -14612 29843 -14556 29877
rect -14522 29843 -14466 29877
rect -14432 29843 -14376 29877
rect -14342 29843 -14286 29877
rect -14252 29843 -14196 29877
rect -14162 29843 -14106 29877
rect -14072 29843 -14016 29877
rect -13982 29843 -13926 29877
rect -13892 29843 -13836 29877
rect -13802 29843 -13628 29877
rect -13594 29843 -13538 29877
rect -13504 29843 -13448 29877
rect -13414 29843 -13358 29877
rect -13324 29843 -13268 29877
rect -13234 29843 -13178 29877
rect -13144 29843 -13088 29877
rect -13054 29843 -12998 29877
rect -12964 29843 -12908 29877
rect -12874 29843 -12818 29877
rect -12784 29843 -12728 29877
rect -12694 29843 -12638 29877
rect -12604 29843 -12548 29877
rect -12514 29843 -12340 29877
rect -12306 29843 -12250 29877
rect -12216 29843 -12160 29877
rect -12126 29843 -12070 29877
rect -12036 29843 -11980 29877
rect -11946 29843 -11890 29877
rect -11856 29843 -11800 29877
rect -11766 29843 -11710 29877
rect -11676 29843 -11620 29877
rect -11586 29843 -11530 29877
rect -11496 29843 -11440 29877
rect -11406 29843 -11350 29877
rect -11316 29843 -11260 29877
rect -11226 29843 -11052 29877
rect -11018 29843 -10962 29877
rect -10928 29843 -10872 29877
rect -10838 29843 -10782 29877
rect -10748 29843 -10692 29877
rect -10658 29843 -10602 29877
rect -10568 29843 -10512 29877
rect -10478 29843 -10422 29877
rect -10388 29843 -10332 29877
rect -10298 29843 -10242 29877
rect -10208 29843 -10152 29877
rect -10118 29843 -10062 29877
rect -10028 29843 -9972 29877
rect -9938 29843 -9764 29877
rect -9730 29843 -9674 29877
rect -9640 29843 -9584 29877
rect -9550 29843 -9494 29877
rect -9460 29843 -9404 29877
rect -9370 29843 -9314 29877
rect -9280 29843 -9224 29877
rect -9190 29843 -9134 29877
rect -9100 29843 -9044 29877
rect -9010 29843 -8954 29877
rect -8920 29843 -8864 29877
rect -8830 29843 -8774 29877
rect -8740 29843 -8684 29877
rect -8650 29843 -8476 29877
rect -8442 29843 -8386 29877
rect -8352 29843 -8296 29877
rect -8262 29843 -8206 29877
rect -8172 29843 -8116 29877
rect -8082 29843 -8026 29877
rect -7992 29843 -7936 29877
rect -7902 29843 -7846 29877
rect -7812 29843 -7756 29877
rect -7722 29843 -7666 29877
rect -7632 29843 -7576 29877
rect -7542 29843 -7486 29877
rect -7452 29843 -7396 29877
rect -7362 29843 -7188 29877
rect -7154 29843 -7098 29877
rect -7064 29843 -7008 29877
rect -6974 29843 -6918 29877
rect -6884 29843 -6828 29877
rect -6794 29843 -6738 29877
rect -6704 29843 -6648 29877
rect -6614 29843 -6558 29877
rect -6524 29843 -6468 29877
rect -6434 29843 -6378 29877
rect -6344 29843 -6288 29877
rect -6254 29843 -6198 29877
rect -6164 29843 -6108 29877
rect -6074 29843 -5900 29877
rect -5866 29843 -5810 29877
rect -5776 29843 -5720 29877
rect -5686 29843 -5630 29877
rect -5596 29843 -5540 29877
rect -5506 29843 -5450 29877
rect -5416 29843 -5360 29877
rect -5326 29843 -5270 29877
rect -5236 29843 -5180 29877
rect -5146 29843 -5090 29877
rect -5056 29843 -5000 29877
rect -4966 29843 -4910 29877
rect -4876 29843 -4820 29877
rect -4786 29843 -4612 29877
rect -4578 29843 -4522 29877
rect -4488 29843 -4432 29877
rect -4398 29843 -4342 29877
rect -4308 29843 -4252 29877
rect -4218 29843 -4162 29877
rect -4128 29843 -4072 29877
rect -4038 29843 -4014 29877
rect -18824 29820 -4014 29843
rect -18824 29809 -4002 29820
rect -18824 29808 -18665 29809
rect -18824 29794 -18722 29808
rect -18824 29760 -18792 29794
rect -18756 29784 -18722 29794
rect -17579 29784 -17377 29809
rect -16291 29784 -16089 29809
rect -15003 29784 -14873 29809
rect -13787 29784 -13585 29809
rect -12499 29784 -12297 29809
rect -11211 29784 -11009 29809
rect -9923 29784 -9721 29809
rect -8635 29784 -8433 29809
rect -7347 29784 -7145 29809
rect -6059 29784 -5857 29809
rect -4771 29784 -4569 29809
rect -18756 29760 -18723 29784
rect -18824 29704 -18723 29760
rect -18824 29670 -18791 29704
rect -18757 29670 -18723 29704
rect -18824 29614 -18723 29670
rect -4128 29704 -4002 29809
rect -4128 29670 -4069 29704
rect -4035 29670 -4002 29704
rect -4128 29661 -4002 29670
rect -18824 29580 -18791 29614
rect -18757 29580 -18723 29614
rect -18824 29524 -18723 29580
rect -18824 29490 -18791 29524
rect -18757 29490 -18723 29524
rect -18824 29434 -18723 29490
rect -18824 29400 -18791 29434
rect -18757 29400 -18723 29434
rect -18824 29344 -18723 29400
rect -18824 29310 -18791 29344
rect -18757 29310 -18723 29344
rect -18824 29254 -18723 29310
rect -18824 29220 -18791 29254
rect -18757 29220 -18723 29254
rect -18824 29164 -18723 29220
rect -18824 29130 -18791 29164
rect -18757 29130 -18723 29164
rect -18824 29074 -18723 29130
rect -18824 29040 -18791 29074
rect -18757 29040 -18723 29074
rect -18824 28984 -18723 29040
rect -18824 28950 -18791 28984
rect -18757 28950 -18723 28984
rect -18824 28894 -18723 28950
rect -18824 28860 -18791 28894
rect -18757 28860 -18723 28894
rect -18824 28804 -18723 28860
rect -18824 28770 -18791 28804
rect -18757 28770 -18723 28804
rect -18824 28723 -18723 28770
rect -4103 29614 -4002 29661
rect -4103 29580 -4069 29614
rect -4035 29580 -4002 29614
rect -4103 29524 -4002 29580
rect -4103 29490 -4069 29524
rect -4035 29490 -4002 29524
rect -4103 29434 -4002 29490
rect -4103 29400 -4069 29434
rect -4035 29400 -4002 29434
rect -4103 29344 -4002 29400
rect -4103 29310 -4069 29344
rect -4035 29310 -4002 29344
rect -4103 29254 -4002 29310
rect -4103 29220 -4069 29254
rect -4035 29220 -4002 29254
rect -4103 29164 -4002 29220
rect -4103 29130 -4069 29164
rect -4035 29130 -4002 29164
rect -4103 29074 -4002 29130
rect -4103 29040 -4069 29074
rect -4035 29040 -4002 29074
rect -4103 28984 -4002 29040
rect -4103 28950 -4069 28984
rect -4035 28950 -4002 28984
rect -4103 28894 -4002 28950
rect -4103 28860 -4069 28894
rect -4035 28860 -4002 28894
rect -4103 28804 -4002 28860
rect -4103 28770 -4069 28804
rect -4035 28770 -4002 28804
rect -18824 28714 -18698 28723
rect -18824 28680 -18791 28714
rect -18757 28680 -18698 28714
rect -18824 28521 -18698 28680
rect -4103 28714 -4002 28770
rect -4103 28680 -4069 28714
rect -4035 28680 -4002 28714
rect -4103 28624 -4002 28680
rect -4103 28590 -4069 28624
rect -4035 28590 -4002 28624
rect -4103 28575 -4002 28590
rect -18824 28506 -18723 28521
rect -18824 28472 -18791 28506
rect -18757 28472 -18723 28506
rect -18824 28416 -18723 28472
rect -18824 28382 -18791 28416
rect -18757 28382 -18723 28416
rect -18824 28326 -18723 28382
rect -4128 28416 -4002 28575
rect -4128 28382 -4069 28416
rect -4035 28382 -4002 28416
rect -4128 28373 -4002 28382
rect -18824 28292 -18791 28326
rect -18757 28292 -18723 28326
rect -18824 28236 -18723 28292
rect -18824 28202 -18791 28236
rect -18757 28202 -18723 28236
rect -18824 28146 -18723 28202
rect -18824 28112 -18791 28146
rect -18757 28112 -18723 28146
rect -18824 28056 -18723 28112
rect -18824 28022 -18791 28056
rect -18757 28022 -18723 28056
rect -18824 27966 -18723 28022
rect -18824 27932 -18791 27966
rect -18757 27932 -18723 27966
rect -18824 27876 -18723 27932
rect -18824 27842 -18791 27876
rect -18757 27842 -18723 27876
rect -18824 27786 -18723 27842
rect -18824 27752 -18791 27786
rect -18757 27752 -18723 27786
rect -18824 27696 -18723 27752
rect -18824 27662 -18791 27696
rect -18757 27662 -18723 27696
rect -18824 27606 -18723 27662
rect -18824 27572 -18791 27606
rect -18757 27572 -18723 27606
rect -18824 27516 -18723 27572
rect -18824 27482 -18791 27516
rect -18757 27482 -18723 27516
rect -18824 27435 -18723 27482
rect -4103 28326 -4002 28373
rect -4103 28292 -4069 28326
rect -4035 28292 -4002 28326
rect -4103 28236 -4002 28292
rect -4103 28202 -4069 28236
rect -4035 28202 -4002 28236
rect -4103 28146 -4002 28202
rect -4103 28112 -4069 28146
rect -4035 28112 -4002 28146
rect -4103 28056 -4002 28112
rect -4103 28022 -4069 28056
rect -4035 28022 -4002 28056
rect -4103 27966 -4002 28022
rect -4103 27932 -4069 27966
rect -4035 27932 -4002 27966
rect -4103 27876 -4002 27932
rect -4103 27842 -4069 27876
rect -4035 27842 -4002 27876
rect -4103 27786 -4002 27842
rect -4103 27752 -4069 27786
rect -4035 27752 -4002 27786
rect -4103 27696 -4002 27752
rect -4103 27662 -4069 27696
rect -4035 27662 -4002 27696
rect -4103 27606 -4002 27662
rect -4103 27572 -4069 27606
rect -4035 27572 -4002 27606
rect -4103 27516 -4002 27572
rect -4103 27482 -4069 27516
rect -4035 27482 -4002 27516
rect -18824 27426 -18698 27435
rect -18824 27392 -18791 27426
rect -18757 27392 -18698 27426
rect -18824 27233 -18698 27392
rect -4103 27426 -4002 27482
rect -4103 27392 -4069 27426
rect -4035 27392 -4002 27426
rect -4103 27336 -4002 27392
rect -4103 27302 -4069 27336
rect -4035 27302 -4002 27336
rect -4103 27287 -4002 27302
rect -18824 27218 -18723 27233
rect -18824 27184 -18791 27218
rect -18757 27184 -18723 27218
rect -18824 27128 -18723 27184
rect -18824 27094 -18791 27128
rect -18757 27094 -18723 27128
rect -18824 27038 -18723 27094
rect -4128 27128 -4002 27287
rect -4128 27094 -4069 27128
rect -4035 27094 -4002 27128
rect -4128 27085 -4002 27094
rect -18824 27004 -18791 27038
rect -18757 27004 -18723 27038
rect -18824 26948 -18723 27004
rect -18824 26914 -18791 26948
rect -18757 26914 -18723 26948
rect -18824 26858 -18723 26914
rect -18824 26824 -18791 26858
rect -18757 26824 -18723 26858
rect -18824 26768 -18723 26824
rect -18824 26734 -18791 26768
rect -18757 26734 -18723 26768
rect -18824 26678 -18723 26734
rect -18824 26644 -18791 26678
rect -18757 26644 -18723 26678
rect -18824 26588 -18723 26644
rect -18824 26554 -18791 26588
rect -18757 26554 -18723 26588
rect -18824 26498 -18723 26554
rect -18824 26464 -18791 26498
rect -18757 26464 -18723 26498
rect -18824 26408 -18723 26464
rect -18824 26374 -18791 26408
rect -18757 26374 -18723 26408
rect -18824 26318 -18723 26374
rect -18824 26284 -18791 26318
rect -18757 26284 -18723 26318
rect -18824 26228 -18723 26284
rect -18824 26194 -18791 26228
rect -18757 26194 -18723 26228
rect -18824 26147 -18723 26194
rect -4103 27038 -4002 27085
rect -4103 27004 -4069 27038
rect -4035 27004 -4002 27038
rect -4103 26948 -4002 27004
rect -4103 26914 -4069 26948
rect -4035 26914 -4002 26948
rect -4103 26858 -4002 26914
rect -4103 26824 -4069 26858
rect -4035 26824 -4002 26858
rect -4103 26768 -4002 26824
rect -4103 26734 -4069 26768
rect -4035 26734 -4002 26768
rect -4103 26678 -4002 26734
rect -4103 26644 -4069 26678
rect -4035 26644 -4002 26678
rect -4103 26588 -4002 26644
rect -4103 26554 -4069 26588
rect -4035 26554 -4002 26588
rect -4103 26498 -4002 26554
rect -4103 26464 -4069 26498
rect -4035 26464 -4002 26498
rect -4103 26408 -4002 26464
rect -4103 26374 -4069 26408
rect -4035 26374 -4002 26408
rect -4103 26318 -4002 26374
rect -4103 26284 -4069 26318
rect -4035 26284 -4002 26318
rect -4103 26228 -4002 26284
rect -4103 26194 -4069 26228
rect -4035 26194 -4002 26228
rect -18824 26138 -18698 26147
rect -18824 26104 -18791 26138
rect -18757 26104 -18698 26138
rect -18824 25945 -18698 26104
rect -4103 26138 -4002 26194
rect -4103 26104 -4069 26138
rect -4035 26104 -4002 26138
rect -4103 26048 -4002 26104
rect -4103 26014 -4069 26048
rect -4035 26014 -4002 26048
rect -4103 25999 -4002 26014
rect -18824 25930 -18723 25945
rect -18824 25896 -18791 25930
rect -18757 25896 -18723 25930
rect -18824 25840 -18723 25896
rect -4128 25912 -4002 25999
rect -4128 25878 -4069 25912
rect -4035 25878 -4002 25912
rect -4128 25869 -4002 25878
rect -18824 25806 -18791 25840
rect -18757 25806 -18723 25840
rect -18824 25750 -18723 25806
rect -18824 25716 -18791 25750
rect -18757 25716 -18723 25750
rect -18824 25660 -18723 25716
rect -18824 25626 -18791 25660
rect -18757 25626 -18723 25660
rect -18824 25570 -18723 25626
rect -18824 25536 -18791 25570
rect -18757 25536 -18723 25570
rect -18824 25480 -18723 25536
rect -18824 25446 -18791 25480
rect -18757 25446 -18723 25480
rect -18824 25390 -18723 25446
rect -18824 25356 -18791 25390
rect -18757 25356 -18723 25390
rect -18824 25300 -18723 25356
rect -18824 25266 -18791 25300
rect -18757 25266 -18723 25300
rect -18824 25210 -18723 25266
rect -18824 25176 -18791 25210
rect -18757 25176 -18723 25210
rect -18824 25120 -18723 25176
rect -18824 25086 -18791 25120
rect -18757 25086 -18723 25120
rect -18824 25030 -18723 25086
rect -18824 24996 -18791 25030
rect -18757 24996 -18723 25030
rect -18824 24940 -18723 24996
rect -18824 24906 -18791 24940
rect -18757 24906 -18723 24940
rect -18824 24859 -18723 24906
rect -4103 25822 -4002 25869
rect -4103 25788 -4069 25822
rect -4035 25788 -4002 25822
rect -4103 25732 -4002 25788
rect -4103 25698 -4069 25732
rect -4035 25698 -4002 25732
rect -4103 25642 -4002 25698
rect -4103 25608 -4069 25642
rect -4035 25608 -4002 25642
rect -4103 25552 -4002 25608
rect -4103 25518 -4069 25552
rect -4035 25518 -4002 25552
rect -4103 25462 -4002 25518
rect -4103 25428 -4069 25462
rect -4035 25428 -4002 25462
rect -4103 25372 -4002 25428
rect -4103 25338 -4069 25372
rect -4035 25338 -4002 25372
rect -4103 25282 -4002 25338
rect -4103 25248 -4069 25282
rect -4035 25248 -4002 25282
rect -4103 25192 -4002 25248
rect -4103 25158 -4069 25192
rect -4035 25158 -4002 25192
rect -4103 25102 -4002 25158
rect -4103 25068 -4069 25102
rect -4035 25068 -4002 25102
rect -4103 25012 -4002 25068
rect -4103 24978 -4069 25012
rect -4035 24978 -4002 25012
rect -4103 24922 -4002 24978
rect -4103 24888 -4069 24922
rect -4035 24888 -4002 24922
rect -18824 24850 -18698 24859
rect -18824 24816 -18791 24850
rect -18757 24816 -18698 24850
rect -18824 24657 -18698 24816
rect -4103 24832 -4002 24888
rect -4103 24798 -4069 24832
rect -4035 24798 -4002 24832
rect -4103 24783 -4002 24798
rect -18824 24642 -18723 24657
rect -18824 24608 -18791 24642
rect -18757 24608 -18723 24642
rect -18824 24552 -18723 24608
rect -4128 24624 -4002 24783
rect -4128 24590 -4069 24624
rect -4035 24590 -4002 24624
rect -4128 24581 -4002 24590
rect -18824 24518 -18791 24552
rect -18757 24518 -18723 24552
rect -18824 24462 -18723 24518
rect -18824 24428 -18791 24462
rect -18757 24428 -18723 24462
rect -18824 24372 -18723 24428
rect -18824 24338 -18791 24372
rect -18757 24338 -18723 24372
rect -18824 24282 -18723 24338
rect -18824 24248 -18791 24282
rect -18757 24248 -18723 24282
rect -18824 24192 -18723 24248
rect -18824 24158 -18791 24192
rect -18757 24158 -18723 24192
rect -18824 24102 -18723 24158
rect -18824 24068 -18791 24102
rect -18757 24068 -18723 24102
rect -18824 24012 -18723 24068
rect -18824 23978 -18791 24012
rect -18757 23978 -18723 24012
rect -18824 23922 -18723 23978
rect -18824 23888 -18791 23922
rect -18757 23888 -18723 23922
rect -18824 23832 -18723 23888
rect -18824 23798 -18791 23832
rect -18757 23798 -18723 23832
rect -18824 23742 -18723 23798
rect -18824 23708 -18791 23742
rect -18757 23708 -18723 23742
rect -18824 23652 -18723 23708
rect -18824 23618 -18791 23652
rect -18757 23618 -18723 23652
rect -18824 23571 -18723 23618
rect -4103 24534 -4002 24581
rect -4103 24500 -4069 24534
rect -4035 24500 -4002 24534
rect -4103 24444 -4002 24500
rect -4103 24410 -4069 24444
rect -4035 24410 -4002 24444
rect -4103 24354 -4002 24410
rect -4103 24320 -4069 24354
rect -4035 24320 -4002 24354
rect -4103 24264 -4002 24320
rect -4103 24230 -4069 24264
rect -4035 24230 -4002 24264
rect -4103 24174 -4002 24230
rect -4103 24140 -4069 24174
rect -4035 24140 -4002 24174
rect -4103 24084 -4002 24140
rect -4103 24050 -4069 24084
rect -4035 24050 -4002 24084
rect -4103 23994 -4002 24050
rect -4103 23960 -4069 23994
rect -4035 23960 -4002 23994
rect -4103 23904 -4002 23960
rect -4103 23870 -4069 23904
rect -4035 23870 -4002 23904
rect -4103 23814 -4002 23870
rect -4103 23780 -4069 23814
rect -4035 23780 -4002 23814
rect -4103 23724 -4002 23780
rect -4103 23690 -4069 23724
rect -4035 23690 -4002 23724
rect -4103 23634 -4002 23690
rect -4103 23600 -4069 23634
rect -4035 23600 -4002 23634
rect -18824 23562 -18698 23571
rect -18824 23528 -18791 23562
rect -18757 23528 -18698 23562
rect -18824 23369 -18698 23528
rect -4103 23544 -4002 23600
rect -4103 23510 -4069 23544
rect -4035 23510 -4002 23544
rect -4103 23495 -4002 23510
rect -18824 23354 -18723 23369
rect -18824 23320 -18791 23354
rect -18757 23320 -18723 23354
rect -18824 23264 -18723 23320
rect -4128 23336 -4002 23495
rect -4128 23302 -4069 23336
rect -4035 23302 -4002 23336
rect -4128 23293 -4002 23302
rect -18824 23230 -18791 23264
rect -18757 23230 -18723 23264
rect -18824 23174 -18723 23230
rect -18824 23140 -18791 23174
rect -18757 23140 -18723 23174
rect -18824 23084 -18723 23140
rect -18824 23050 -18791 23084
rect -18757 23050 -18723 23084
rect -18824 22994 -18723 23050
rect -18824 22960 -18791 22994
rect -18757 22960 -18723 22994
rect -18824 22904 -18723 22960
rect -18824 22870 -18791 22904
rect -18757 22870 -18723 22904
rect -18824 22814 -18723 22870
rect -18824 22780 -18791 22814
rect -18757 22780 -18723 22814
rect -18824 22724 -18723 22780
rect -18824 22690 -18791 22724
rect -18757 22690 -18723 22724
rect -18824 22634 -18723 22690
rect -18824 22600 -18791 22634
rect -18757 22600 -18723 22634
rect -18824 22544 -18723 22600
rect -18824 22510 -18791 22544
rect -18757 22510 -18723 22544
rect -18824 22454 -18723 22510
rect -18824 22420 -18791 22454
rect -18757 22420 -18723 22454
rect -18824 22364 -18723 22420
rect -18824 22330 -18791 22364
rect -18757 22330 -18723 22364
rect -18824 22283 -18723 22330
rect -4103 23246 -4002 23293
rect -4103 23212 -4069 23246
rect -4035 23212 -4002 23246
rect -4103 23156 -4002 23212
rect -4103 23122 -4069 23156
rect -4035 23122 -4002 23156
rect -4103 23066 -4002 23122
rect -4103 23032 -4069 23066
rect -4035 23032 -4002 23066
rect -4103 22976 -4002 23032
rect -4103 22942 -4069 22976
rect -4035 22942 -4002 22976
rect -4103 22886 -4002 22942
rect -4103 22852 -4069 22886
rect -4035 22852 -4002 22886
rect -4103 22796 -4002 22852
rect -4103 22762 -4069 22796
rect -4035 22762 -4002 22796
rect -4103 22706 -4002 22762
rect -4103 22672 -4069 22706
rect -4035 22672 -4002 22706
rect -4103 22616 -4002 22672
rect -4103 22582 -4069 22616
rect -4035 22582 -4002 22616
rect -4103 22526 -4002 22582
rect -4103 22492 -4069 22526
rect -4035 22492 -4002 22526
rect -4103 22436 -4002 22492
rect -4103 22402 -4069 22436
rect -4035 22402 -4002 22436
rect -4103 22346 -4002 22402
rect -4103 22312 -4069 22346
rect -4035 22312 -4002 22346
rect -18824 22274 -18698 22283
rect -18824 22240 -18791 22274
rect -18757 22240 -18698 22274
rect -18824 22081 -18698 22240
rect -4103 22256 -4002 22312
rect -4103 22222 -4069 22256
rect -4035 22222 -4002 22256
rect -4103 22207 -4002 22222
rect -18824 22066 -18723 22081
rect -18824 22032 -18791 22066
rect -18757 22032 -18723 22066
rect -18824 21976 -18723 22032
rect -4128 22048 -4002 22207
rect -4128 22014 -4069 22048
rect -4035 22014 -4002 22048
rect -4128 22005 -4002 22014
rect -18824 21942 -18791 21976
rect -18757 21942 -18723 21976
rect -18824 21886 -18723 21942
rect -18824 21852 -18791 21886
rect -18757 21852 -18723 21886
rect -18824 21796 -18723 21852
rect -18824 21762 -18791 21796
rect -18757 21762 -18723 21796
rect -18824 21706 -18723 21762
rect -18824 21672 -18791 21706
rect -18757 21672 -18723 21706
rect -18824 21616 -18723 21672
rect -18824 21582 -18791 21616
rect -18757 21582 -18723 21616
rect -18824 21526 -18723 21582
rect -18824 21492 -18791 21526
rect -18757 21492 -18723 21526
rect -18824 21436 -18723 21492
rect -18824 21402 -18791 21436
rect -18757 21402 -18723 21436
rect -18824 21346 -18723 21402
rect -18824 21312 -18791 21346
rect -18757 21312 -18723 21346
rect -18824 21256 -18723 21312
rect -18824 21222 -18791 21256
rect -18757 21222 -18723 21256
rect -18824 21166 -18723 21222
rect -18824 21132 -18791 21166
rect -18757 21132 -18723 21166
rect -18824 21076 -18723 21132
rect -18824 21042 -18791 21076
rect -18757 21042 -18723 21076
rect -18824 20995 -18723 21042
rect -4103 21958 -4002 22005
rect -4103 21924 -4069 21958
rect -4035 21924 -4002 21958
rect -4103 21868 -4002 21924
rect -4103 21834 -4069 21868
rect -4035 21834 -4002 21868
rect -4103 21778 -4002 21834
rect -4103 21744 -4069 21778
rect -4035 21744 -4002 21778
rect -4103 21688 -4002 21744
rect -4103 21654 -4069 21688
rect -4035 21654 -4002 21688
rect -4103 21598 -4002 21654
rect -4103 21564 -4069 21598
rect -4035 21564 -4002 21598
rect -4103 21508 -4002 21564
rect -4103 21474 -4069 21508
rect -4035 21474 -4002 21508
rect -4103 21418 -4002 21474
rect -4103 21384 -4069 21418
rect -4035 21384 -4002 21418
rect -4103 21328 -4002 21384
rect -4103 21294 -4069 21328
rect -4035 21294 -4002 21328
rect -4103 21238 -4002 21294
rect -4103 21204 -4069 21238
rect -4035 21204 -4002 21238
rect -4103 21148 -4002 21204
rect -4103 21114 -4069 21148
rect -4035 21114 -4002 21148
rect -4103 21058 -4002 21114
rect -4103 21024 -4069 21058
rect -4035 21024 -4002 21058
rect -18824 20986 -18698 20995
rect -18824 20952 -18791 20986
rect -18757 20952 -18698 20986
rect -18824 20793 -18698 20952
rect -4103 20968 -4002 21024
rect -4103 20934 -4069 20968
rect -4035 20934 -4002 20968
rect -4103 20919 -4002 20934
rect -18824 20778 -18723 20793
rect -18824 20744 -18791 20778
rect -18757 20744 -18723 20778
rect -18824 20688 -18723 20744
rect -4128 20760 -4002 20919
rect -4128 20726 -4069 20760
rect -4035 20726 -4002 20760
rect -4128 20717 -4002 20726
rect -18824 20654 -18791 20688
rect -18757 20654 -18723 20688
rect -18824 20598 -18723 20654
rect -18824 20564 -18791 20598
rect -18757 20564 -18723 20598
rect -18824 20508 -18723 20564
rect -18824 20474 -18791 20508
rect -18757 20474 -18723 20508
rect -18824 20418 -18723 20474
rect -18824 20384 -18791 20418
rect -18757 20384 -18723 20418
rect -18824 20328 -18723 20384
rect -18824 20294 -18791 20328
rect -18757 20294 -18723 20328
rect -18824 20238 -18723 20294
rect -18824 20204 -18791 20238
rect -18757 20204 -18723 20238
rect -18824 20148 -18723 20204
rect -18824 20114 -18791 20148
rect -18757 20114 -18723 20148
rect -18824 20058 -18723 20114
rect -18824 20024 -18791 20058
rect -18757 20024 -18723 20058
rect -18824 19968 -18723 20024
rect -18824 19934 -18791 19968
rect -18757 19934 -18723 19968
rect -18824 19878 -18723 19934
rect -18824 19844 -18791 19878
rect -18757 19844 -18723 19878
rect -18824 19788 -18723 19844
rect -18824 19754 -18791 19788
rect -18757 19754 -18723 19788
rect -18824 19707 -18723 19754
rect -4103 20670 -4002 20717
rect -4103 20636 -4069 20670
rect -4035 20636 -4002 20670
rect -4103 20580 -4002 20636
rect -4103 20546 -4069 20580
rect -4035 20546 -4002 20580
rect -4103 20490 -4002 20546
rect -4103 20456 -4069 20490
rect -4035 20456 -4002 20490
rect -4103 20400 -4002 20456
rect -4103 20366 -4069 20400
rect -4035 20366 -4002 20400
rect -4103 20310 -4002 20366
rect -4103 20276 -4069 20310
rect -4035 20276 -4002 20310
rect -4103 20220 -4002 20276
rect -4103 20186 -4069 20220
rect -4035 20186 -4002 20220
rect -4103 20130 -4002 20186
rect -4103 20096 -4069 20130
rect -4035 20096 -4002 20130
rect -4103 20040 -4002 20096
rect -4103 20006 -4069 20040
rect -4035 20006 -4002 20040
rect -4103 19950 -4002 20006
rect -4103 19916 -4069 19950
rect -4035 19916 -4002 19950
rect -4103 19860 -4002 19916
rect -4103 19826 -4069 19860
rect -4035 19826 -4002 19860
rect -4103 19770 -4002 19826
rect -4103 19736 -4069 19770
rect -4035 19736 -4002 19770
rect -18824 19698 -18698 19707
rect -18824 19664 -18791 19698
rect -18757 19664 -18698 19698
rect -18824 19505 -18698 19664
rect -4103 19680 -4002 19736
rect -4103 19646 -4069 19680
rect -4035 19646 -4002 19680
rect -4103 19631 -4002 19646
rect -18824 19490 -18723 19505
rect -18824 19456 -18791 19490
rect -18757 19456 -18723 19490
rect -18824 19400 -18723 19456
rect -4128 19472 -4002 19631
rect -4128 19438 -4069 19472
rect -4035 19438 -4002 19472
rect -4128 19429 -4002 19438
rect -18824 19366 -18791 19400
rect -18757 19366 -18723 19400
rect -18824 19310 -18723 19366
rect -18824 19276 -18791 19310
rect -18757 19276 -18723 19310
rect -18824 19220 -18723 19276
rect -18824 19186 -18791 19220
rect -18757 19186 -18723 19220
rect -18824 19130 -18723 19186
rect -18824 19096 -18791 19130
rect -18757 19096 -18723 19130
rect -18824 19040 -18723 19096
rect -18824 19006 -18791 19040
rect -18757 19006 -18723 19040
rect -18824 18950 -18723 19006
rect -18824 18916 -18791 18950
rect -18757 18916 -18723 18950
rect -18824 18860 -18723 18916
rect -18824 18826 -18791 18860
rect -18757 18826 -18723 18860
rect -18824 18770 -18723 18826
rect -18824 18736 -18791 18770
rect -18757 18736 -18723 18770
rect -18824 18680 -18723 18736
rect -18824 18646 -18791 18680
rect -18757 18646 -18723 18680
rect -18824 18590 -18723 18646
rect -18824 18556 -18791 18590
rect -18757 18556 -18723 18590
rect -18824 18500 -18723 18556
rect -18824 18466 -18791 18500
rect -18757 18466 -18723 18500
rect -18824 18419 -18723 18466
rect -4103 19382 -4002 19429
rect -4103 19348 -4069 19382
rect -4035 19348 -4002 19382
rect -4103 19292 -4002 19348
rect -4103 19258 -4069 19292
rect -4035 19258 -4002 19292
rect -4103 19202 -4002 19258
rect -4103 19168 -4069 19202
rect -4035 19168 -4002 19202
rect -4103 19112 -4002 19168
rect -4103 19078 -4069 19112
rect -4035 19078 -4002 19112
rect -4103 19022 -4002 19078
rect -4103 18988 -4069 19022
rect -4035 18988 -4002 19022
rect -4103 18932 -4002 18988
rect -4103 18898 -4069 18932
rect -4035 18898 -4002 18932
rect -4103 18842 -4002 18898
rect -4103 18808 -4069 18842
rect -4035 18808 -4002 18842
rect -4103 18752 -4002 18808
rect -4103 18718 -4069 18752
rect -4035 18718 -4002 18752
rect -4103 18662 -4002 18718
rect -4103 18628 -4069 18662
rect -4035 18628 -4002 18662
rect -4103 18572 -4002 18628
rect -4103 18538 -4069 18572
rect -4035 18538 -4002 18572
rect -4103 18482 -4002 18538
rect -4103 18448 -4069 18482
rect -4035 18448 -4002 18482
rect -18824 18410 -18698 18419
rect -18824 18376 -18791 18410
rect -18757 18376 -18698 18410
rect -18824 18217 -18698 18376
rect -4103 18392 -4002 18448
rect -4103 18358 -4069 18392
rect -4035 18358 -4002 18392
rect -4103 18343 -4002 18358
rect -18824 18202 -18723 18217
rect -18824 18168 -18791 18202
rect -18757 18168 -18723 18202
rect -18824 18112 -18723 18168
rect -4128 18184 -4002 18343
rect -4128 18150 -4069 18184
rect -4035 18150 -4002 18184
rect -4128 18141 -4002 18150
rect -18824 18078 -18791 18112
rect -18757 18078 -18723 18112
rect -18824 18022 -18723 18078
rect -18824 17988 -18791 18022
rect -18757 17988 -18723 18022
rect -18824 17932 -18723 17988
rect -18824 17898 -18791 17932
rect -18757 17898 -18723 17932
rect -18824 17842 -18723 17898
rect -18824 17808 -18791 17842
rect -18757 17808 -18723 17842
rect -18824 17752 -18723 17808
rect -18824 17718 -18791 17752
rect -18757 17718 -18723 17752
rect -18824 17662 -18723 17718
rect -18824 17628 -18791 17662
rect -18757 17628 -18723 17662
rect -18824 17572 -18723 17628
rect -18824 17538 -18791 17572
rect -18757 17538 -18723 17572
rect -18824 17482 -18723 17538
rect -18824 17448 -18791 17482
rect -18757 17448 -18723 17482
rect -18824 17392 -18723 17448
rect -18824 17358 -18791 17392
rect -18757 17358 -18723 17392
rect -18824 17302 -18723 17358
rect -18824 17268 -18791 17302
rect -18757 17268 -18723 17302
rect -18824 17212 -18723 17268
rect -18824 17178 -18791 17212
rect -18757 17178 -18723 17212
rect -18824 17131 -18723 17178
rect -4103 18094 -4002 18141
rect -4103 18060 -4069 18094
rect -4035 18060 -4002 18094
rect -4103 18004 -4002 18060
rect -4103 17970 -4069 18004
rect -4035 17970 -4002 18004
rect -4103 17914 -4002 17970
rect -4103 17880 -4069 17914
rect -4035 17880 -4002 17914
rect -4103 17824 -4002 17880
rect -4103 17790 -4069 17824
rect -4035 17790 -4002 17824
rect -4103 17734 -4002 17790
rect -4103 17700 -4069 17734
rect -4035 17700 -4002 17734
rect -4103 17644 -4002 17700
rect -4103 17610 -4069 17644
rect -4035 17610 -4002 17644
rect -4103 17554 -4002 17610
rect -4103 17520 -4069 17554
rect -4035 17520 -4002 17554
rect -4103 17464 -4002 17520
rect -4103 17430 -4069 17464
rect -4035 17430 -4002 17464
rect -4103 17374 -4002 17430
rect -4103 17340 -4069 17374
rect -4035 17340 -4002 17374
rect -4103 17284 -4002 17340
rect -4103 17250 -4069 17284
rect -4035 17250 -4002 17284
rect -4103 17194 -4002 17250
rect -4103 17160 -4069 17194
rect -4035 17160 -4002 17194
rect -18824 17122 -18698 17131
rect -18824 17088 -18791 17122
rect -18757 17088 -18698 17122
rect -18824 17001 -18698 17088
rect -4103 17104 -4002 17160
rect -4103 17070 -4069 17104
rect -4035 17070 -4002 17104
rect -4103 17055 -4002 17070
rect -18824 16986 -18723 17001
rect -18824 16952 -18791 16986
rect -18757 16952 -18723 16986
rect -18824 16896 -18723 16952
rect -18824 16862 -18791 16896
rect -18757 16862 -18723 16896
rect -18824 16806 -18723 16862
rect -4128 16896 -4002 17055
rect -4128 16862 -4069 16896
rect -4035 16862 -4002 16896
rect -4128 16853 -4002 16862
rect -18824 16772 -18791 16806
rect -18757 16772 -18723 16806
rect -18824 16716 -18723 16772
rect -18824 16682 -18791 16716
rect -18757 16682 -18723 16716
rect -18824 16626 -18723 16682
rect -18824 16592 -18791 16626
rect -18757 16592 -18723 16626
rect -18824 16536 -18723 16592
rect -18824 16502 -18791 16536
rect -18757 16502 -18723 16536
rect -18824 16446 -18723 16502
rect -18824 16412 -18791 16446
rect -18757 16412 -18723 16446
rect -18824 16356 -18723 16412
rect -18824 16322 -18791 16356
rect -18757 16322 -18723 16356
rect -18824 16266 -18723 16322
rect -18824 16232 -18791 16266
rect -18757 16232 -18723 16266
rect -18824 16176 -18723 16232
rect -18824 16142 -18791 16176
rect -18757 16142 -18723 16176
rect -18824 16086 -18723 16142
rect -18824 16052 -18791 16086
rect -18757 16052 -18723 16086
rect -18824 15996 -18723 16052
rect -18824 15962 -18791 15996
rect -18757 15962 -18723 15996
rect -18824 15915 -18723 15962
rect -4103 16806 -4002 16853
rect -4103 16772 -4069 16806
rect -4035 16772 -4002 16806
rect -4103 16716 -4002 16772
rect -4103 16682 -4069 16716
rect -4035 16682 -4002 16716
rect -4103 16626 -4002 16682
rect -4103 16592 -4069 16626
rect -4035 16592 -4002 16626
rect -4103 16536 -4002 16592
rect -4103 16502 -4069 16536
rect -4035 16502 -4002 16536
rect -4103 16446 -4002 16502
rect -4103 16412 -4069 16446
rect -4035 16412 -4002 16446
rect -4103 16356 -4002 16412
rect -4103 16322 -4069 16356
rect -4035 16322 -4002 16356
rect -4103 16266 -4002 16322
rect -4103 16232 -4069 16266
rect -4035 16232 -4002 16266
rect -4103 16176 -4002 16232
rect -4103 16142 -4069 16176
rect -4035 16142 -4002 16176
rect -4103 16086 -4002 16142
rect -4103 16052 -4069 16086
rect -4035 16052 -4002 16086
rect -4103 15996 -4002 16052
rect -4103 15962 -4069 15996
rect -4035 15962 -4002 15996
rect -18824 15906 -18698 15915
rect -18824 15872 -18791 15906
rect -18757 15872 -18698 15906
rect -18824 15713 -18698 15872
rect -4103 15906 -4002 15962
rect -4103 15872 -4069 15906
rect -4035 15872 -4002 15906
rect -4103 15816 -4002 15872
rect -4103 15782 -4069 15816
rect -4035 15782 -4002 15816
rect -4103 15767 -4002 15782
rect -18824 15698 -18723 15713
rect -18824 15664 -18791 15698
rect -18757 15664 -18723 15698
rect -18824 15608 -18723 15664
rect -18824 15574 -18791 15608
rect -18757 15574 -18723 15608
rect -18824 15518 -18723 15574
rect -4128 15608 -4002 15767
rect -4128 15574 -4069 15608
rect -4035 15574 -4002 15608
rect -4128 15565 -4002 15574
rect -18824 15484 -18791 15518
rect -18757 15484 -18723 15518
rect -18824 15428 -18723 15484
rect -18824 15394 -18791 15428
rect -18757 15394 -18723 15428
rect -18824 15338 -18723 15394
rect -18824 15304 -18791 15338
rect -18757 15304 -18723 15338
rect -18824 15248 -18723 15304
rect -18824 15214 -18791 15248
rect -18757 15214 -18723 15248
rect -18824 15158 -18723 15214
rect -18824 15124 -18791 15158
rect -18757 15124 -18723 15158
rect -18824 15068 -18723 15124
rect -18824 15034 -18791 15068
rect -18757 15034 -18723 15068
rect -18824 14978 -18723 15034
rect -18824 14944 -18791 14978
rect -18757 14944 -18723 14978
rect -18824 14888 -18723 14944
rect -18824 14854 -18791 14888
rect -18757 14854 -18723 14888
rect -18824 14798 -18723 14854
rect -18824 14764 -18791 14798
rect -18757 14764 -18723 14798
rect -18824 14708 -18723 14764
rect -18824 14674 -18791 14708
rect -18757 14674 -18723 14708
rect -18824 14627 -18723 14674
rect -4103 15518 -4002 15565
rect -4103 15484 -4069 15518
rect -4035 15484 -4002 15518
rect -4103 15428 -4002 15484
rect -4103 15394 -4069 15428
rect -4035 15394 -4002 15428
rect -4103 15338 -4002 15394
rect -4103 15304 -4069 15338
rect -4035 15304 -4002 15338
rect -4103 15248 -4002 15304
rect -4103 15214 -4069 15248
rect -4035 15214 -4002 15248
rect -4103 15158 -4002 15214
rect -4103 15124 -4069 15158
rect -4035 15124 -4002 15158
rect -4103 15068 -4002 15124
rect -4103 15034 -4069 15068
rect -4035 15034 -4002 15068
rect -4103 14978 -4002 15034
rect -4103 14944 -4069 14978
rect -4035 14944 -4002 14978
rect -4103 14888 -4002 14944
rect -4103 14854 -4069 14888
rect -4035 14854 -4002 14888
rect -4103 14798 -4002 14854
rect -4103 14764 -4069 14798
rect -4035 14764 -4002 14798
rect -4103 14708 -4002 14764
rect -4103 14674 -4069 14708
rect -4035 14674 -4002 14708
rect -18824 14618 -18698 14627
rect -18824 14584 -18791 14618
rect -18757 14584 -18698 14618
rect -18824 14425 -18698 14584
rect -4103 14618 -4002 14674
rect -4103 14584 -4069 14618
rect -4035 14584 -4002 14618
rect -4103 14528 -4002 14584
rect -4103 14494 -4069 14528
rect -4035 14494 -4002 14528
rect -4103 14479 -4002 14494
rect -18824 14410 -18723 14425
rect -18824 14376 -18791 14410
rect -18757 14376 -18723 14410
rect -18824 14320 -18723 14376
rect -18824 14286 -18791 14320
rect -18757 14286 -18723 14320
rect -18824 14230 -18723 14286
rect -4128 14320 -4002 14479
rect -4128 14286 -4069 14320
rect -4035 14286 -4002 14320
rect -4128 14277 -4002 14286
rect -18824 14196 -18791 14230
rect -18757 14196 -18723 14230
rect -18824 14140 -18723 14196
rect -18824 14106 -18791 14140
rect -18757 14106 -18723 14140
rect -18824 14050 -18723 14106
rect -18824 14016 -18791 14050
rect -18757 14016 -18723 14050
rect -18824 13960 -18723 14016
rect -18824 13926 -18791 13960
rect -18757 13926 -18723 13960
rect -18824 13870 -18723 13926
rect -18824 13836 -18791 13870
rect -18757 13836 -18723 13870
rect -18824 13780 -18723 13836
rect -18824 13746 -18791 13780
rect -18757 13746 -18723 13780
rect -18824 13690 -18723 13746
rect -18824 13656 -18791 13690
rect -18757 13656 -18723 13690
rect -18824 13600 -18723 13656
rect -18824 13566 -18791 13600
rect -18757 13566 -18723 13600
rect -18824 13510 -18723 13566
rect -18824 13476 -18791 13510
rect -18757 13476 -18723 13510
rect -18824 13420 -18723 13476
rect -18824 13386 -18791 13420
rect -18757 13386 -18723 13420
rect -18824 13339 -18723 13386
rect -4103 14230 -4002 14277
rect -4103 14196 -4069 14230
rect -4035 14196 -4002 14230
rect -4103 14140 -4002 14196
rect -4103 14106 -4069 14140
rect -4035 14106 -4002 14140
rect -4103 14050 -4002 14106
rect -4103 14016 -4069 14050
rect -4035 14016 -4002 14050
rect -4103 13960 -4002 14016
rect -4103 13926 -4069 13960
rect -4035 13926 -4002 13960
rect -4103 13870 -4002 13926
rect -4103 13836 -4069 13870
rect -4035 13836 -4002 13870
rect -4103 13780 -4002 13836
rect -4103 13746 -4069 13780
rect -4035 13746 -4002 13780
rect -4103 13690 -4002 13746
rect -4103 13656 -4069 13690
rect -4035 13656 -4002 13690
rect -4103 13600 -4002 13656
rect -4103 13566 -4069 13600
rect -4035 13566 -4002 13600
rect -4103 13510 -4002 13566
rect -4103 13476 -4069 13510
rect -4035 13476 -4002 13510
rect -4103 13420 -4002 13476
rect -4103 13386 -4069 13420
rect -4035 13386 -4002 13420
rect -18824 13330 -18698 13339
rect -18824 13296 -18791 13330
rect -18757 13296 -18698 13330
rect -18824 13191 -18698 13296
rect -4103 13330 -4002 13386
rect -4103 13296 -4069 13330
rect -4035 13296 -4002 13330
rect -4103 13240 -4002 13296
rect -4103 13216 -4070 13240
rect -18257 13191 -18055 13216
rect -16969 13191 -16767 13216
rect -15681 13191 -15479 13216
rect -14393 13191 -14191 13216
rect -13105 13191 -12903 13216
rect -11817 13191 -11615 13216
rect -10529 13191 -10327 13216
rect -9241 13191 -9039 13216
rect -7953 13191 -7823 13216
rect -6737 13191 -6535 13216
rect -5449 13191 -5247 13216
rect -4104 13206 -4070 13216
rect -4034 13206 -4002 13240
rect -4104 13192 -4002 13206
rect -4161 13191 -4002 13192
rect -18824 13180 -4002 13191
rect -18812 13157 -4002 13180
rect -18812 13123 -18788 13157
rect -18754 13123 -18698 13157
rect -18664 13123 -18608 13157
rect -18574 13123 -18518 13157
rect -18484 13123 -18428 13157
rect -18394 13123 -18338 13157
rect -18304 13123 -18248 13157
rect -18214 13123 -18040 13157
rect -18006 13123 -17950 13157
rect -17916 13123 -17860 13157
rect -17826 13123 -17770 13157
rect -17736 13123 -17680 13157
rect -17646 13123 -17590 13157
rect -17556 13123 -17500 13157
rect -17466 13123 -17410 13157
rect -17376 13123 -17320 13157
rect -17286 13123 -17230 13157
rect -17196 13123 -17140 13157
rect -17106 13123 -17050 13157
rect -17016 13123 -16960 13157
rect -16926 13123 -16752 13157
rect -16718 13123 -16662 13157
rect -16628 13123 -16572 13157
rect -16538 13123 -16482 13157
rect -16448 13123 -16392 13157
rect -16358 13123 -16302 13157
rect -16268 13123 -16212 13157
rect -16178 13123 -16122 13157
rect -16088 13123 -16032 13157
rect -15998 13123 -15942 13157
rect -15908 13123 -15852 13157
rect -15818 13123 -15762 13157
rect -15728 13123 -15672 13157
rect -15638 13123 -15464 13157
rect -15430 13123 -15374 13157
rect -15340 13123 -15284 13157
rect -15250 13123 -15194 13157
rect -15160 13123 -15104 13157
rect -15070 13123 -15014 13157
rect -14980 13123 -14924 13157
rect -14890 13123 -14834 13157
rect -14800 13123 -14744 13157
rect -14710 13123 -14654 13157
rect -14620 13123 -14564 13157
rect -14530 13123 -14474 13157
rect -14440 13123 -14384 13157
rect -14350 13123 -14176 13157
rect -14142 13123 -14086 13157
rect -14052 13123 -13996 13157
rect -13962 13123 -13906 13157
rect -13872 13123 -13816 13157
rect -13782 13123 -13726 13157
rect -13692 13123 -13636 13157
rect -13602 13123 -13546 13157
rect -13512 13123 -13456 13157
rect -13422 13123 -13366 13157
rect -13332 13123 -13276 13157
rect -13242 13123 -13186 13157
rect -13152 13123 -13096 13157
rect -13062 13123 -12888 13157
rect -12854 13123 -12798 13157
rect -12764 13123 -12708 13157
rect -12674 13123 -12618 13157
rect -12584 13123 -12528 13157
rect -12494 13123 -12438 13157
rect -12404 13123 -12348 13157
rect -12314 13123 -12258 13157
rect -12224 13123 -12168 13157
rect -12134 13123 -12078 13157
rect -12044 13123 -11988 13157
rect -11954 13123 -11898 13157
rect -11864 13123 -11808 13157
rect -11774 13123 -11600 13157
rect -11566 13123 -11510 13157
rect -11476 13123 -11420 13157
rect -11386 13123 -11330 13157
rect -11296 13123 -11240 13157
rect -11206 13123 -11150 13157
rect -11116 13123 -11060 13157
rect -11026 13123 -10970 13157
rect -10936 13123 -10880 13157
rect -10846 13123 -10790 13157
rect -10756 13123 -10700 13157
rect -10666 13123 -10610 13157
rect -10576 13123 -10520 13157
rect -10486 13123 -10312 13157
rect -10278 13123 -10222 13157
rect -10188 13123 -10132 13157
rect -10098 13123 -10042 13157
rect -10008 13123 -9952 13157
rect -9918 13123 -9862 13157
rect -9828 13123 -9772 13157
rect -9738 13123 -9682 13157
rect -9648 13123 -9592 13157
rect -9558 13123 -9502 13157
rect -9468 13123 -9412 13157
rect -9378 13123 -9322 13157
rect -9288 13123 -9232 13157
rect -9198 13123 -9024 13157
rect -8990 13123 -8934 13157
rect -8900 13123 -8844 13157
rect -8810 13123 -8754 13157
rect -8720 13123 -8664 13157
rect -8630 13123 -8574 13157
rect -8540 13123 -8484 13157
rect -8450 13123 -8394 13157
rect -8360 13123 -8304 13157
rect -8270 13123 -8214 13157
rect -8180 13123 -8124 13157
rect -8090 13123 -8034 13157
rect -8000 13123 -7944 13157
rect -7910 13123 -7808 13157
rect -7774 13123 -7718 13157
rect -7684 13123 -7628 13157
rect -7594 13123 -7538 13157
rect -7504 13123 -7448 13157
rect -7414 13123 -7358 13157
rect -7324 13123 -7268 13157
rect -7234 13123 -7178 13157
rect -7144 13123 -7088 13157
rect -7054 13123 -6998 13157
rect -6964 13123 -6908 13157
rect -6874 13123 -6818 13157
rect -6784 13123 -6728 13157
rect -6694 13123 -6520 13157
rect -6486 13123 -6430 13157
rect -6396 13123 -6340 13157
rect -6306 13123 -6250 13157
rect -6216 13123 -6160 13157
rect -6126 13123 -6070 13157
rect -6036 13123 -5980 13157
rect -5946 13123 -5890 13157
rect -5856 13123 -5800 13157
rect -5766 13123 -5710 13157
rect -5676 13123 -5620 13157
rect -5586 13123 -5530 13157
rect -5496 13123 -5440 13157
rect -5406 13123 -5232 13157
rect -5198 13123 -5142 13157
rect -5108 13123 -5052 13157
rect -5018 13123 -4962 13157
rect -4928 13123 -4872 13157
rect -4838 13123 -4782 13157
rect -4748 13123 -4692 13157
rect -4658 13123 -4602 13157
rect -4568 13123 -4512 13157
rect -4478 13123 -4422 13157
rect -4388 13123 -4332 13157
rect -4298 13123 -4242 13157
rect -4208 13123 -4152 13157
rect -4118 13123 -4002 13157
rect -18812 13090 -4002 13123
rect -18812 13084 -18766 13090
<< psubdiffcont >>
rect -18708 29843 -18674 29877
rect -18618 29843 -18584 29877
rect -18528 29843 -18494 29877
rect -18438 29843 -18404 29877
rect -18348 29843 -18314 29877
rect -18258 29843 -18224 29877
rect -18168 29843 -18134 29877
rect -18078 29843 -18044 29877
rect -17988 29843 -17954 29877
rect -17898 29843 -17864 29877
rect -17808 29843 -17774 29877
rect -17718 29843 -17684 29877
rect -17628 29843 -17594 29877
rect -17420 29843 -17386 29877
rect -17330 29843 -17296 29877
rect -17240 29843 -17206 29877
rect -17150 29843 -17116 29877
rect -17060 29843 -17026 29877
rect -16970 29843 -16936 29877
rect -16880 29843 -16846 29877
rect -16790 29843 -16756 29877
rect -16700 29843 -16666 29877
rect -16610 29843 -16576 29877
rect -16520 29843 -16486 29877
rect -16430 29843 -16396 29877
rect -16340 29843 -16306 29877
rect -16132 29843 -16098 29877
rect -16042 29843 -16008 29877
rect -15952 29843 -15918 29877
rect -15862 29843 -15828 29877
rect -15772 29843 -15738 29877
rect -15682 29843 -15648 29877
rect -15592 29843 -15558 29877
rect -15502 29843 -15468 29877
rect -15412 29843 -15378 29877
rect -15322 29843 -15288 29877
rect -15232 29843 -15198 29877
rect -15142 29843 -15108 29877
rect -15052 29843 -15018 29877
rect -14916 29843 -14882 29877
rect -14826 29843 -14792 29877
rect -14736 29843 -14702 29877
rect -14646 29843 -14612 29877
rect -14556 29843 -14522 29877
rect -14466 29843 -14432 29877
rect -14376 29843 -14342 29877
rect -14286 29843 -14252 29877
rect -14196 29843 -14162 29877
rect -14106 29843 -14072 29877
rect -14016 29843 -13982 29877
rect -13926 29843 -13892 29877
rect -13836 29843 -13802 29877
rect -13628 29843 -13594 29877
rect -13538 29843 -13504 29877
rect -13448 29843 -13414 29877
rect -13358 29843 -13324 29877
rect -13268 29843 -13234 29877
rect -13178 29843 -13144 29877
rect -13088 29843 -13054 29877
rect -12998 29843 -12964 29877
rect -12908 29843 -12874 29877
rect -12818 29843 -12784 29877
rect -12728 29843 -12694 29877
rect -12638 29843 -12604 29877
rect -12548 29843 -12514 29877
rect -12340 29843 -12306 29877
rect -12250 29843 -12216 29877
rect -12160 29843 -12126 29877
rect -12070 29843 -12036 29877
rect -11980 29843 -11946 29877
rect -11890 29843 -11856 29877
rect -11800 29843 -11766 29877
rect -11710 29843 -11676 29877
rect -11620 29843 -11586 29877
rect -11530 29843 -11496 29877
rect -11440 29843 -11406 29877
rect -11350 29843 -11316 29877
rect -11260 29843 -11226 29877
rect -11052 29843 -11018 29877
rect -10962 29843 -10928 29877
rect -10872 29843 -10838 29877
rect -10782 29843 -10748 29877
rect -10692 29843 -10658 29877
rect -10602 29843 -10568 29877
rect -10512 29843 -10478 29877
rect -10422 29843 -10388 29877
rect -10332 29843 -10298 29877
rect -10242 29843 -10208 29877
rect -10152 29843 -10118 29877
rect -10062 29843 -10028 29877
rect -9972 29843 -9938 29877
rect -9764 29843 -9730 29877
rect -9674 29843 -9640 29877
rect -9584 29843 -9550 29877
rect -9494 29843 -9460 29877
rect -9404 29843 -9370 29877
rect -9314 29843 -9280 29877
rect -9224 29843 -9190 29877
rect -9134 29843 -9100 29877
rect -9044 29843 -9010 29877
rect -8954 29843 -8920 29877
rect -8864 29843 -8830 29877
rect -8774 29843 -8740 29877
rect -8684 29843 -8650 29877
rect -8476 29843 -8442 29877
rect -8386 29843 -8352 29877
rect -8296 29843 -8262 29877
rect -8206 29843 -8172 29877
rect -8116 29843 -8082 29877
rect -8026 29843 -7992 29877
rect -7936 29843 -7902 29877
rect -7846 29843 -7812 29877
rect -7756 29843 -7722 29877
rect -7666 29843 -7632 29877
rect -7576 29843 -7542 29877
rect -7486 29843 -7452 29877
rect -7396 29843 -7362 29877
rect -7188 29843 -7154 29877
rect -7098 29843 -7064 29877
rect -7008 29843 -6974 29877
rect -6918 29843 -6884 29877
rect -6828 29843 -6794 29877
rect -6738 29843 -6704 29877
rect -6648 29843 -6614 29877
rect -6558 29843 -6524 29877
rect -6468 29843 -6434 29877
rect -6378 29843 -6344 29877
rect -6288 29843 -6254 29877
rect -6198 29843 -6164 29877
rect -6108 29843 -6074 29877
rect -5900 29843 -5866 29877
rect -5810 29843 -5776 29877
rect -5720 29843 -5686 29877
rect -5630 29843 -5596 29877
rect -5540 29843 -5506 29877
rect -5450 29843 -5416 29877
rect -5360 29843 -5326 29877
rect -5270 29843 -5236 29877
rect -5180 29843 -5146 29877
rect -5090 29843 -5056 29877
rect -5000 29843 -4966 29877
rect -4910 29843 -4876 29877
rect -4820 29843 -4786 29877
rect -4612 29843 -4578 29877
rect -4522 29843 -4488 29877
rect -4432 29843 -4398 29877
rect -4342 29843 -4308 29877
rect -4252 29843 -4218 29877
rect -4162 29843 -4128 29877
rect -4072 29843 -4038 29877
rect -18792 29760 -18756 29794
rect -18791 29670 -18757 29704
rect -4069 29670 -4035 29704
rect -18791 29580 -18757 29614
rect -18791 29490 -18757 29524
rect -18791 29400 -18757 29434
rect -18791 29310 -18757 29344
rect -18791 29220 -18757 29254
rect -18791 29130 -18757 29164
rect -18791 29040 -18757 29074
rect -18791 28950 -18757 28984
rect -18791 28860 -18757 28894
rect -18791 28770 -18757 28804
rect -4069 29580 -4035 29614
rect -4069 29490 -4035 29524
rect -4069 29400 -4035 29434
rect -4069 29310 -4035 29344
rect -4069 29220 -4035 29254
rect -4069 29130 -4035 29164
rect -4069 29040 -4035 29074
rect -4069 28950 -4035 28984
rect -4069 28860 -4035 28894
rect -4069 28770 -4035 28804
rect -18791 28680 -18757 28714
rect -4069 28680 -4035 28714
rect -4069 28590 -4035 28624
rect -18791 28472 -18757 28506
rect -18791 28382 -18757 28416
rect -4069 28382 -4035 28416
rect -18791 28292 -18757 28326
rect -18791 28202 -18757 28236
rect -18791 28112 -18757 28146
rect -18791 28022 -18757 28056
rect -18791 27932 -18757 27966
rect -18791 27842 -18757 27876
rect -18791 27752 -18757 27786
rect -18791 27662 -18757 27696
rect -18791 27572 -18757 27606
rect -18791 27482 -18757 27516
rect -4069 28292 -4035 28326
rect -4069 28202 -4035 28236
rect -4069 28112 -4035 28146
rect -4069 28022 -4035 28056
rect -4069 27932 -4035 27966
rect -4069 27842 -4035 27876
rect -4069 27752 -4035 27786
rect -4069 27662 -4035 27696
rect -4069 27572 -4035 27606
rect -4069 27482 -4035 27516
rect -18791 27392 -18757 27426
rect -4069 27392 -4035 27426
rect -4069 27302 -4035 27336
rect -18791 27184 -18757 27218
rect -18791 27094 -18757 27128
rect -4069 27094 -4035 27128
rect -18791 27004 -18757 27038
rect -18791 26914 -18757 26948
rect -18791 26824 -18757 26858
rect -18791 26734 -18757 26768
rect -18791 26644 -18757 26678
rect -18791 26554 -18757 26588
rect -18791 26464 -18757 26498
rect -18791 26374 -18757 26408
rect -18791 26284 -18757 26318
rect -18791 26194 -18757 26228
rect -4069 27004 -4035 27038
rect -4069 26914 -4035 26948
rect -4069 26824 -4035 26858
rect -4069 26734 -4035 26768
rect -4069 26644 -4035 26678
rect -4069 26554 -4035 26588
rect -4069 26464 -4035 26498
rect -4069 26374 -4035 26408
rect -4069 26284 -4035 26318
rect -4069 26194 -4035 26228
rect -18791 26104 -18757 26138
rect -4069 26104 -4035 26138
rect -4069 26014 -4035 26048
rect -18791 25896 -18757 25930
rect -4069 25878 -4035 25912
rect -18791 25806 -18757 25840
rect -18791 25716 -18757 25750
rect -18791 25626 -18757 25660
rect -18791 25536 -18757 25570
rect -18791 25446 -18757 25480
rect -18791 25356 -18757 25390
rect -18791 25266 -18757 25300
rect -18791 25176 -18757 25210
rect -18791 25086 -18757 25120
rect -18791 24996 -18757 25030
rect -18791 24906 -18757 24940
rect -4069 25788 -4035 25822
rect -4069 25698 -4035 25732
rect -4069 25608 -4035 25642
rect -4069 25518 -4035 25552
rect -4069 25428 -4035 25462
rect -4069 25338 -4035 25372
rect -4069 25248 -4035 25282
rect -4069 25158 -4035 25192
rect -4069 25068 -4035 25102
rect -4069 24978 -4035 25012
rect -4069 24888 -4035 24922
rect -18791 24816 -18757 24850
rect -4069 24798 -4035 24832
rect -18791 24608 -18757 24642
rect -4069 24590 -4035 24624
rect -18791 24518 -18757 24552
rect -18791 24428 -18757 24462
rect -18791 24338 -18757 24372
rect -18791 24248 -18757 24282
rect -18791 24158 -18757 24192
rect -18791 24068 -18757 24102
rect -18791 23978 -18757 24012
rect -18791 23888 -18757 23922
rect -18791 23798 -18757 23832
rect -18791 23708 -18757 23742
rect -18791 23618 -18757 23652
rect -4069 24500 -4035 24534
rect -4069 24410 -4035 24444
rect -4069 24320 -4035 24354
rect -4069 24230 -4035 24264
rect -4069 24140 -4035 24174
rect -4069 24050 -4035 24084
rect -4069 23960 -4035 23994
rect -4069 23870 -4035 23904
rect -4069 23780 -4035 23814
rect -4069 23690 -4035 23724
rect -4069 23600 -4035 23634
rect -18791 23528 -18757 23562
rect -4069 23510 -4035 23544
rect -18791 23320 -18757 23354
rect -4069 23302 -4035 23336
rect -18791 23230 -18757 23264
rect -18791 23140 -18757 23174
rect -18791 23050 -18757 23084
rect -18791 22960 -18757 22994
rect -18791 22870 -18757 22904
rect -18791 22780 -18757 22814
rect -18791 22690 -18757 22724
rect -18791 22600 -18757 22634
rect -18791 22510 -18757 22544
rect -18791 22420 -18757 22454
rect -18791 22330 -18757 22364
rect -4069 23212 -4035 23246
rect -4069 23122 -4035 23156
rect -4069 23032 -4035 23066
rect -4069 22942 -4035 22976
rect -4069 22852 -4035 22886
rect -4069 22762 -4035 22796
rect -4069 22672 -4035 22706
rect -4069 22582 -4035 22616
rect -4069 22492 -4035 22526
rect -4069 22402 -4035 22436
rect -4069 22312 -4035 22346
rect -18791 22240 -18757 22274
rect -4069 22222 -4035 22256
rect -18791 22032 -18757 22066
rect -4069 22014 -4035 22048
rect -18791 21942 -18757 21976
rect -18791 21852 -18757 21886
rect -18791 21762 -18757 21796
rect -18791 21672 -18757 21706
rect -18791 21582 -18757 21616
rect -18791 21492 -18757 21526
rect -18791 21402 -18757 21436
rect -18791 21312 -18757 21346
rect -18791 21222 -18757 21256
rect -18791 21132 -18757 21166
rect -18791 21042 -18757 21076
rect -4069 21924 -4035 21958
rect -4069 21834 -4035 21868
rect -4069 21744 -4035 21778
rect -4069 21654 -4035 21688
rect -4069 21564 -4035 21598
rect -4069 21474 -4035 21508
rect -4069 21384 -4035 21418
rect -4069 21294 -4035 21328
rect -4069 21204 -4035 21238
rect -4069 21114 -4035 21148
rect -4069 21024 -4035 21058
rect -18791 20952 -18757 20986
rect -4069 20934 -4035 20968
rect -18791 20744 -18757 20778
rect -4069 20726 -4035 20760
rect -18791 20654 -18757 20688
rect -18791 20564 -18757 20598
rect -18791 20474 -18757 20508
rect -18791 20384 -18757 20418
rect -18791 20294 -18757 20328
rect -18791 20204 -18757 20238
rect -18791 20114 -18757 20148
rect -18791 20024 -18757 20058
rect -18791 19934 -18757 19968
rect -18791 19844 -18757 19878
rect -18791 19754 -18757 19788
rect -4069 20636 -4035 20670
rect -4069 20546 -4035 20580
rect -4069 20456 -4035 20490
rect -4069 20366 -4035 20400
rect -4069 20276 -4035 20310
rect -4069 20186 -4035 20220
rect -4069 20096 -4035 20130
rect -4069 20006 -4035 20040
rect -4069 19916 -4035 19950
rect -4069 19826 -4035 19860
rect -4069 19736 -4035 19770
rect -18791 19664 -18757 19698
rect -4069 19646 -4035 19680
rect -18791 19456 -18757 19490
rect -4069 19438 -4035 19472
rect -18791 19366 -18757 19400
rect -18791 19276 -18757 19310
rect -18791 19186 -18757 19220
rect -18791 19096 -18757 19130
rect -18791 19006 -18757 19040
rect -18791 18916 -18757 18950
rect -18791 18826 -18757 18860
rect -18791 18736 -18757 18770
rect -18791 18646 -18757 18680
rect -18791 18556 -18757 18590
rect -18791 18466 -18757 18500
rect -4069 19348 -4035 19382
rect -4069 19258 -4035 19292
rect -4069 19168 -4035 19202
rect -4069 19078 -4035 19112
rect -4069 18988 -4035 19022
rect -4069 18898 -4035 18932
rect -4069 18808 -4035 18842
rect -4069 18718 -4035 18752
rect -4069 18628 -4035 18662
rect -4069 18538 -4035 18572
rect -4069 18448 -4035 18482
rect -18791 18376 -18757 18410
rect -4069 18358 -4035 18392
rect -18791 18168 -18757 18202
rect -4069 18150 -4035 18184
rect -18791 18078 -18757 18112
rect -18791 17988 -18757 18022
rect -18791 17898 -18757 17932
rect -18791 17808 -18757 17842
rect -18791 17718 -18757 17752
rect -18791 17628 -18757 17662
rect -18791 17538 -18757 17572
rect -18791 17448 -18757 17482
rect -18791 17358 -18757 17392
rect -18791 17268 -18757 17302
rect -18791 17178 -18757 17212
rect -4069 18060 -4035 18094
rect -4069 17970 -4035 18004
rect -4069 17880 -4035 17914
rect -4069 17790 -4035 17824
rect -4069 17700 -4035 17734
rect -4069 17610 -4035 17644
rect -4069 17520 -4035 17554
rect -4069 17430 -4035 17464
rect -4069 17340 -4035 17374
rect -4069 17250 -4035 17284
rect -4069 17160 -4035 17194
rect -18791 17088 -18757 17122
rect -4069 17070 -4035 17104
rect -18791 16952 -18757 16986
rect -18791 16862 -18757 16896
rect -4069 16862 -4035 16896
rect -18791 16772 -18757 16806
rect -18791 16682 -18757 16716
rect -18791 16592 -18757 16626
rect -18791 16502 -18757 16536
rect -18791 16412 -18757 16446
rect -18791 16322 -18757 16356
rect -18791 16232 -18757 16266
rect -18791 16142 -18757 16176
rect -18791 16052 -18757 16086
rect -18791 15962 -18757 15996
rect -4069 16772 -4035 16806
rect -4069 16682 -4035 16716
rect -4069 16592 -4035 16626
rect -4069 16502 -4035 16536
rect -4069 16412 -4035 16446
rect -4069 16322 -4035 16356
rect -4069 16232 -4035 16266
rect -4069 16142 -4035 16176
rect -4069 16052 -4035 16086
rect -4069 15962 -4035 15996
rect -18791 15872 -18757 15906
rect -4069 15872 -4035 15906
rect -4069 15782 -4035 15816
rect -18791 15664 -18757 15698
rect -18791 15574 -18757 15608
rect -4069 15574 -4035 15608
rect -18791 15484 -18757 15518
rect -18791 15394 -18757 15428
rect -18791 15304 -18757 15338
rect -18791 15214 -18757 15248
rect -18791 15124 -18757 15158
rect -18791 15034 -18757 15068
rect -18791 14944 -18757 14978
rect -18791 14854 -18757 14888
rect -18791 14764 -18757 14798
rect -18791 14674 -18757 14708
rect -4069 15484 -4035 15518
rect -4069 15394 -4035 15428
rect -4069 15304 -4035 15338
rect -4069 15214 -4035 15248
rect -4069 15124 -4035 15158
rect -4069 15034 -4035 15068
rect -4069 14944 -4035 14978
rect -4069 14854 -4035 14888
rect -4069 14764 -4035 14798
rect -4069 14674 -4035 14708
rect -18791 14584 -18757 14618
rect -4069 14584 -4035 14618
rect -4069 14494 -4035 14528
rect -18791 14376 -18757 14410
rect -18791 14286 -18757 14320
rect -4069 14286 -4035 14320
rect -18791 14196 -18757 14230
rect -18791 14106 -18757 14140
rect -18791 14016 -18757 14050
rect -18791 13926 -18757 13960
rect -18791 13836 -18757 13870
rect -18791 13746 -18757 13780
rect -18791 13656 -18757 13690
rect -18791 13566 -18757 13600
rect -18791 13476 -18757 13510
rect -18791 13386 -18757 13420
rect -4069 14196 -4035 14230
rect -4069 14106 -4035 14140
rect -4069 14016 -4035 14050
rect -4069 13926 -4035 13960
rect -4069 13836 -4035 13870
rect -4069 13746 -4035 13780
rect -4069 13656 -4035 13690
rect -4069 13566 -4035 13600
rect -4069 13476 -4035 13510
rect -4069 13386 -4035 13420
rect -18791 13296 -18757 13330
rect -4069 13296 -4035 13330
rect -4070 13206 -4034 13240
rect -18788 13123 -18754 13157
rect -18698 13123 -18664 13157
rect -18608 13123 -18574 13157
rect -18518 13123 -18484 13157
rect -18428 13123 -18394 13157
rect -18338 13123 -18304 13157
rect -18248 13123 -18214 13157
rect -18040 13123 -18006 13157
rect -17950 13123 -17916 13157
rect -17860 13123 -17826 13157
rect -17770 13123 -17736 13157
rect -17680 13123 -17646 13157
rect -17590 13123 -17556 13157
rect -17500 13123 -17466 13157
rect -17410 13123 -17376 13157
rect -17320 13123 -17286 13157
rect -17230 13123 -17196 13157
rect -17140 13123 -17106 13157
rect -17050 13123 -17016 13157
rect -16960 13123 -16926 13157
rect -16752 13123 -16718 13157
rect -16662 13123 -16628 13157
rect -16572 13123 -16538 13157
rect -16482 13123 -16448 13157
rect -16392 13123 -16358 13157
rect -16302 13123 -16268 13157
rect -16212 13123 -16178 13157
rect -16122 13123 -16088 13157
rect -16032 13123 -15998 13157
rect -15942 13123 -15908 13157
rect -15852 13123 -15818 13157
rect -15762 13123 -15728 13157
rect -15672 13123 -15638 13157
rect -15464 13123 -15430 13157
rect -15374 13123 -15340 13157
rect -15284 13123 -15250 13157
rect -15194 13123 -15160 13157
rect -15104 13123 -15070 13157
rect -15014 13123 -14980 13157
rect -14924 13123 -14890 13157
rect -14834 13123 -14800 13157
rect -14744 13123 -14710 13157
rect -14654 13123 -14620 13157
rect -14564 13123 -14530 13157
rect -14474 13123 -14440 13157
rect -14384 13123 -14350 13157
rect -14176 13123 -14142 13157
rect -14086 13123 -14052 13157
rect -13996 13123 -13962 13157
rect -13906 13123 -13872 13157
rect -13816 13123 -13782 13157
rect -13726 13123 -13692 13157
rect -13636 13123 -13602 13157
rect -13546 13123 -13512 13157
rect -13456 13123 -13422 13157
rect -13366 13123 -13332 13157
rect -13276 13123 -13242 13157
rect -13186 13123 -13152 13157
rect -13096 13123 -13062 13157
rect -12888 13123 -12854 13157
rect -12798 13123 -12764 13157
rect -12708 13123 -12674 13157
rect -12618 13123 -12584 13157
rect -12528 13123 -12494 13157
rect -12438 13123 -12404 13157
rect -12348 13123 -12314 13157
rect -12258 13123 -12224 13157
rect -12168 13123 -12134 13157
rect -12078 13123 -12044 13157
rect -11988 13123 -11954 13157
rect -11898 13123 -11864 13157
rect -11808 13123 -11774 13157
rect -11600 13123 -11566 13157
rect -11510 13123 -11476 13157
rect -11420 13123 -11386 13157
rect -11330 13123 -11296 13157
rect -11240 13123 -11206 13157
rect -11150 13123 -11116 13157
rect -11060 13123 -11026 13157
rect -10970 13123 -10936 13157
rect -10880 13123 -10846 13157
rect -10790 13123 -10756 13157
rect -10700 13123 -10666 13157
rect -10610 13123 -10576 13157
rect -10520 13123 -10486 13157
rect -10312 13123 -10278 13157
rect -10222 13123 -10188 13157
rect -10132 13123 -10098 13157
rect -10042 13123 -10008 13157
rect -9952 13123 -9918 13157
rect -9862 13123 -9828 13157
rect -9772 13123 -9738 13157
rect -9682 13123 -9648 13157
rect -9592 13123 -9558 13157
rect -9502 13123 -9468 13157
rect -9412 13123 -9378 13157
rect -9322 13123 -9288 13157
rect -9232 13123 -9198 13157
rect -9024 13123 -8990 13157
rect -8934 13123 -8900 13157
rect -8844 13123 -8810 13157
rect -8754 13123 -8720 13157
rect -8664 13123 -8630 13157
rect -8574 13123 -8540 13157
rect -8484 13123 -8450 13157
rect -8394 13123 -8360 13157
rect -8304 13123 -8270 13157
rect -8214 13123 -8180 13157
rect -8124 13123 -8090 13157
rect -8034 13123 -8000 13157
rect -7944 13123 -7910 13157
rect -7808 13123 -7774 13157
rect -7718 13123 -7684 13157
rect -7628 13123 -7594 13157
rect -7538 13123 -7504 13157
rect -7448 13123 -7414 13157
rect -7358 13123 -7324 13157
rect -7268 13123 -7234 13157
rect -7178 13123 -7144 13157
rect -7088 13123 -7054 13157
rect -6998 13123 -6964 13157
rect -6908 13123 -6874 13157
rect -6818 13123 -6784 13157
rect -6728 13123 -6694 13157
rect -6520 13123 -6486 13157
rect -6430 13123 -6396 13157
rect -6340 13123 -6306 13157
rect -6250 13123 -6216 13157
rect -6160 13123 -6126 13157
rect -6070 13123 -6036 13157
rect -5980 13123 -5946 13157
rect -5890 13123 -5856 13157
rect -5800 13123 -5766 13157
rect -5710 13123 -5676 13157
rect -5620 13123 -5586 13157
rect -5530 13123 -5496 13157
rect -5440 13123 -5406 13157
rect -5232 13123 -5198 13157
rect -5142 13123 -5108 13157
rect -5052 13123 -5018 13157
rect -4962 13123 -4928 13157
rect -4872 13123 -4838 13157
rect -4782 13123 -4748 13157
rect -4692 13123 -4658 13157
rect -4602 13123 -4568 13157
rect -4512 13123 -4478 13157
rect -4422 13123 -4388 13157
rect -4332 13123 -4298 13157
rect -4242 13123 -4208 13157
rect -4152 13123 -4118 13157
<< locali >>
rect -1712 30474 4232 30568
rect -4102 29910 -4002 29916
rect -18824 29877 -4002 29910
rect -18824 29843 -18708 29877
rect -18674 29843 -18618 29877
rect -18584 29843 -18528 29877
rect -18494 29843 -18438 29877
rect -18404 29843 -18348 29877
rect -18314 29843 -18258 29877
rect -18224 29843 -18168 29877
rect -18134 29843 -18078 29877
rect -18044 29843 -17988 29877
rect -17954 29843 -17898 29877
rect -17864 29843 -17808 29877
rect -17774 29843 -17718 29877
rect -17684 29843 -17628 29877
rect -17594 29843 -17420 29877
rect -17386 29843 -17330 29877
rect -17296 29843 -17240 29877
rect -17206 29843 -17150 29877
rect -17116 29843 -17060 29877
rect -17026 29843 -16970 29877
rect -16936 29843 -16880 29877
rect -16846 29843 -16790 29877
rect -16756 29843 -16700 29877
rect -16666 29843 -16610 29877
rect -16576 29843 -16520 29877
rect -16486 29843 -16430 29877
rect -16396 29843 -16340 29877
rect -16306 29843 -16132 29877
rect -16098 29843 -16042 29877
rect -16008 29843 -15952 29877
rect -15918 29843 -15862 29877
rect -15828 29843 -15772 29877
rect -15738 29843 -15682 29877
rect -15648 29843 -15592 29877
rect -15558 29843 -15502 29877
rect -15468 29843 -15412 29877
rect -15378 29843 -15322 29877
rect -15288 29843 -15232 29877
rect -15198 29843 -15142 29877
rect -15108 29843 -15052 29877
rect -15018 29843 -14916 29877
rect -14882 29843 -14826 29877
rect -14792 29843 -14736 29877
rect -14702 29843 -14646 29877
rect -14612 29843 -14556 29877
rect -14522 29843 -14466 29877
rect -14432 29843 -14376 29877
rect -14342 29843 -14286 29877
rect -14252 29843 -14196 29877
rect -14162 29843 -14106 29877
rect -14072 29843 -14016 29877
rect -13982 29843 -13926 29877
rect -13892 29843 -13836 29877
rect -13802 29843 -13628 29877
rect -13594 29843 -13538 29877
rect -13504 29843 -13448 29877
rect -13414 29843 -13358 29877
rect -13324 29843 -13268 29877
rect -13234 29843 -13178 29877
rect -13144 29843 -13088 29877
rect -13054 29843 -12998 29877
rect -12964 29843 -12908 29877
rect -12874 29843 -12818 29877
rect -12784 29843 -12728 29877
rect -12694 29843 -12638 29877
rect -12604 29843 -12548 29877
rect -12514 29843 -12340 29877
rect -12306 29843 -12250 29877
rect -12216 29843 -12160 29877
rect -12126 29843 -12070 29877
rect -12036 29843 -11980 29877
rect -11946 29843 -11890 29877
rect -11856 29843 -11800 29877
rect -11766 29843 -11710 29877
rect -11676 29843 -11620 29877
rect -11586 29843 -11530 29877
rect -11496 29843 -11440 29877
rect -11406 29843 -11350 29877
rect -11316 29843 -11260 29877
rect -11226 29843 -11052 29877
rect -11018 29843 -10962 29877
rect -10928 29843 -10872 29877
rect -10838 29843 -10782 29877
rect -10748 29843 -10692 29877
rect -10658 29843 -10602 29877
rect -10568 29843 -10512 29877
rect -10478 29843 -10422 29877
rect -10388 29843 -10332 29877
rect -10298 29843 -10242 29877
rect -10208 29843 -10152 29877
rect -10118 29843 -10062 29877
rect -10028 29843 -9972 29877
rect -9938 29843 -9764 29877
rect -9730 29843 -9674 29877
rect -9640 29843 -9584 29877
rect -9550 29843 -9494 29877
rect -9460 29843 -9404 29877
rect -9370 29843 -9314 29877
rect -9280 29843 -9224 29877
rect -9190 29843 -9134 29877
rect -9100 29843 -9044 29877
rect -9010 29843 -8954 29877
rect -8920 29843 -8864 29877
rect -8830 29843 -8774 29877
rect -8740 29843 -8684 29877
rect -8650 29843 -8476 29877
rect -8442 29843 -8386 29877
rect -8352 29843 -8296 29877
rect -8262 29843 -8206 29877
rect -8172 29843 -8116 29877
rect -8082 29843 -8026 29877
rect -7992 29843 -7936 29877
rect -7902 29843 -7846 29877
rect -7812 29843 -7756 29877
rect -7722 29843 -7666 29877
rect -7632 29843 -7576 29877
rect -7542 29843 -7486 29877
rect -7452 29843 -7396 29877
rect -7362 29843 -7188 29877
rect -7154 29843 -7098 29877
rect -7064 29843 -7008 29877
rect -6974 29843 -6918 29877
rect -6884 29843 -6828 29877
rect -6794 29843 -6738 29877
rect -6704 29843 -6648 29877
rect -6614 29843 -6558 29877
rect -6524 29843 -6468 29877
rect -6434 29843 -6378 29877
rect -6344 29843 -6288 29877
rect -6254 29843 -6198 29877
rect -6164 29843 -6108 29877
rect -6074 29843 -5900 29877
rect -5866 29843 -5810 29877
rect -5776 29843 -5720 29877
rect -5686 29843 -5630 29877
rect -5596 29843 -5540 29877
rect -5506 29843 -5450 29877
rect -5416 29843 -5360 29877
rect -5326 29843 -5270 29877
rect -5236 29843 -5180 29877
rect -5146 29843 -5090 29877
rect -5056 29843 -5000 29877
rect -4966 29843 -4910 29877
rect -4876 29843 -4820 29877
rect -4786 29843 -4612 29877
rect -4578 29843 -4522 29877
rect -4488 29843 -4432 29877
rect -4398 29843 -4342 29877
rect -4308 29843 -4252 29877
rect -4218 29843 -4162 29877
rect -4128 29843 -4072 29877
rect -4038 29843 -4002 29877
rect -18824 29811 -4002 29843
rect -18824 29808 -18667 29811
rect -18824 29794 -18722 29808
rect -18824 29760 -18792 29794
rect -18756 29784 -18722 29794
rect -17577 29784 -17379 29811
rect -16289 29784 -16091 29811
rect -15001 29784 -14875 29811
rect -13785 29784 -13587 29811
rect -12497 29784 -12299 29811
rect -11209 29784 -11011 29811
rect -9921 29784 -9723 29811
rect -8633 29784 -8435 29811
rect -7345 29784 -7147 29811
rect -6057 29784 -5859 29811
rect -4769 29784 -4571 29811
rect -18756 29760 -18725 29784
rect -18824 29704 -18725 29760
rect -18824 29670 -18791 29704
rect -18757 29670 -18725 29704
rect -18824 29614 -18725 29670
rect -4128 29704 -4002 29811
rect -4128 29670 -4069 29704
rect -4035 29670 -4002 29704
rect -4128 29663 -4002 29670
rect -4102 29658 -4002 29663
rect -18824 29580 -18791 29614
rect -18757 29580 -18725 29614
rect -18824 29524 -18725 29580
rect -18824 29490 -18791 29524
rect -18757 29490 -18725 29524
rect -18824 29434 -18725 29490
rect -18824 29400 -18791 29434
rect -18757 29400 -18725 29434
rect -18824 29344 -18725 29400
rect -18824 29310 -18791 29344
rect -18757 29310 -18725 29344
rect -18824 29254 -18725 29310
rect -18824 29220 -18791 29254
rect -18757 29220 -18725 29254
rect -18824 29164 -18725 29220
rect -18824 29130 -18791 29164
rect -18757 29130 -18725 29164
rect -18824 29074 -18725 29130
rect -18824 29040 -18791 29074
rect -18757 29040 -18725 29074
rect -18824 28984 -18725 29040
rect -18824 28950 -18791 28984
rect -18757 28950 -18725 28984
rect -18824 28894 -18725 28950
rect -18824 28860 -18791 28894
rect -18757 28860 -18725 28894
rect -18824 28804 -18725 28860
rect -18824 28770 -18791 28804
rect -18757 28770 -18725 28804
rect -18824 28721 -18725 28770
rect -4101 29614 -4002 29658
rect -4101 29580 -4069 29614
rect -4035 29580 -4002 29614
rect -4101 29524 -4002 29580
rect -4101 29490 -4069 29524
rect -4035 29490 -4002 29524
rect -4101 29434 -4002 29490
rect -4101 29400 -4069 29434
rect -4035 29400 -4002 29434
rect -4101 29344 -4002 29400
rect -4101 29310 -4069 29344
rect -4035 29310 -4002 29344
rect -4101 29254 -4002 29310
rect -4101 29220 -4069 29254
rect -4035 29220 -4002 29254
rect -4101 29164 -4002 29220
rect -4101 29130 -4069 29164
rect -4035 29130 -4002 29164
rect -4101 29074 -4002 29130
rect -4101 29040 -4069 29074
rect -4035 29040 -4002 29074
rect -4101 28984 -4002 29040
rect -4101 28950 -4069 28984
rect -4035 28950 -4002 28984
rect -4101 28894 -4002 28950
rect -4101 28860 -4069 28894
rect -4035 28860 -4002 28894
rect -4101 28804 -4002 28860
rect -4101 28770 -4069 28804
rect -4035 28770 -4002 28804
rect -18824 28714 -18698 28721
rect -18824 28680 -18791 28714
rect -18757 28680 -18698 28714
rect -18824 28523 -18698 28680
rect -4101 28714 -4002 28770
rect -4101 28680 -4069 28714
rect -4035 28680 -4002 28714
rect -4101 28624 -4002 28680
rect -4101 28590 -4069 28624
rect -4035 28590 -4002 28624
rect -4101 28573 -4002 28590
rect -18824 28506 -18725 28523
rect -18824 28472 -18791 28506
rect -18757 28472 -18725 28506
rect -18824 28416 -18725 28472
rect -18824 28382 -18791 28416
rect -18757 28382 -18725 28416
rect -18824 28326 -18725 28382
rect -4128 28416 -4002 28573
rect -4128 28382 -4069 28416
rect -4035 28382 -4002 28416
rect -4128 28375 -4002 28382
rect -18824 28292 -18791 28326
rect -18757 28292 -18725 28326
rect -18824 28236 -18725 28292
rect -18824 28202 -18791 28236
rect -18757 28202 -18725 28236
rect -18824 28146 -18725 28202
rect -18824 28112 -18791 28146
rect -18757 28112 -18725 28146
rect -18824 28056 -18725 28112
rect -18824 28022 -18791 28056
rect -18757 28022 -18725 28056
rect -18824 27966 -18725 28022
rect -18824 27932 -18791 27966
rect -18757 27932 -18725 27966
rect -18824 27876 -18725 27932
rect -18824 27842 -18791 27876
rect -18757 27842 -18725 27876
rect -18824 27786 -18725 27842
rect -18824 27752 -18791 27786
rect -18757 27752 -18725 27786
rect -18824 27696 -18725 27752
rect -18824 27662 -18791 27696
rect -18757 27662 -18725 27696
rect -18824 27606 -18725 27662
rect -18824 27572 -18791 27606
rect -18757 27572 -18725 27606
rect -18824 27516 -18725 27572
rect -18824 27482 -18791 27516
rect -18757 27482 -18725 27516
rect -18824 27433 -18725 27482
rect -4101 28326 -4002 28375
rect -4101 28292 -4069 28326
rect -4035 28292 -4002 28326
rect -4101 28236 -4002 28292
rect -4101 28202 -4069 28236
rect -4035 28202 -4002 28236
rect -4101 28146 -4002 28202
rect -4101 28112 -4069 28146
rect -4035 28112 -4002 28146
rect -4101 28056 -4002 28112
rect -4101 28022 -4069 28056
rect -4035 28022 -4002 28056
rect -4101 27966 -4002 28022
rect -4101 27932 -4069 27966
rect -4035 27932 -4002 27966
rect -4101 27876 -4002 27932
rect -4101 27842 -4069 27876
rect -4035 27842 -4002 27876
rect -4101 27786 -4002 27842
rect -4101 27752 -4069 27786
rect -4035 27752 -4002 27786
rect -4101 27696 -4002 27752
rect -4101 27662 -4069 27696
rect -4035 27662 -4002 27696
rect -4101 27606 -4002 27662
rect -4101 27572 -4069 27606
rect -4035 27572 -4002 27606
rect -4101 27516 -4002 27572
rect -4101 27482 -4069 27516
rect -4035 27482 -4002 27516
rect -18824 27426 -18698 27433
rect -18824 27392 -18791 27426
rect -18757 27392 -18698 27426
rect -18824 27235 -18698 27392
rect -4101 27426 -4002 27482
rect -4101 27392 -4069 27426
rect -4035 27392 -4002 27426
rect -4101 27336 -4002 27392
rect -4101 27302 -4069 27336
rect -4035 27302 -4002 27336
rect -4101 27285 -4002 27302
rect -18824 27218 -18725 27235
rect -18824 27184 -18791 27218
rect -18757 27184 -18725 27218
rect -18824 27128 -18725 27184
rect -18824 27094 -18791 27128
rect -18757 27094 -18725 27128
rect -18824 27038 -18725 27094
rect -4128 27128 -4002 27285
rect -4128 27094 -4069 27128
rect -4035 27094 -4002 27128
rect -4128 27087 -4002 27094
rect -18824 27004 -18791 27038
rect -18757 27004 -18725 27038
rect -18824 26948 -18725 27004
rect -18824 26914 -18791 26948
rect -18757 26914 -18725 26948
rect -18824 26858 -18725 26914
rect -18824 26824 -18791 26858
rect -18757 26824 -18725 26858
rect -18824 26768 -18725 26824
rect -18824 26734 -18791 26768
rect -18757 26734 -18725 26768
rect -18824 26678 -18725 26734
rect -18824 26644 -18791 26678
rect -18757 26644 -18725 26678
rect -18824 26588 -18725 26644
rect -18824 26554 -18791 26588
rect -18757 26554 -18725 26588
rect -18824 26498 -18725 26554
rect -18824 26464 -18791 26498
rect -18757 26464 -18725 26498
rect -18824 26408 -18725 26464
rect -18824 26374 -18791 26408
rect -18757 26374 -18725 26408
rect -18824 26318 -18725 26374
rect -18824 26284 -18791 26318
rect -18757 26284 -18725 26318
rect -18824 26228 -18725 26284
rect -18824 26194 -18791 26228
rect -18757 26194 -18725 26228
rect -18824 26145 -18725 26194
rect -4101 27038 -4002 27087
rect -4101 27004 -4069 27038
rect -4035 27004 -4002 27038
rect -4101 26948 -4002 27004
rect -4101 26914 -4069 26948
rect -4035 26914 -4002 26948
rect -4101 26858 -4002 26914
rect -4101 26824 -4069 26858
rect -4035 26824 -4002 26858
rect -4101 26768 -4002 26824
rect -4101 26734 -4069 26768
rect -4035 26734 -4002 26768
rect -4101 26678 -4002 26734
rect -4101 26644 -4069 26678
rect -4035 26644 -4002 26678
rect -4101 26588 -4002 26644
rect -4101 26554 -4069 26588
rect -4035 26554 -4002 26588
rect -4101 26498 -4002 26554
rect -4101 26464 -4069 26498
rect -4035 26464 -4002 26498
rect -4101 26408 -4002 26464
rect -4101 26374 -4069 26408
rect -4035 26374 -4002 26408
rect -4101 26318 -4002 26374
rect -4101 26284 -4069 26318
rect -4035 26284 -4002 26318
rect -4101 26228 -4002 26284
rect -4101 26194 -4069 26228
rect -4035 26194 -4002 26228
rect -18824 26138 -18698 26145
rect -18824 26104 -18791 26138
rect -18757 26104 -18698 26138
rect -18824 25947 -18698 26104
rect -4101 26138 -4002 26194
rect -4101 26104 -4069 26138
rect -4035 26104 -4002 26138
rect -4101 26048 -4002 26104
rect -4101 26014 -4069 26048
rect -4035 26014 -4002 26048
rect -4101 25997 -4002 26014
rect -18824 25930 -18725 25947
rect -18824 25896 -18791 25930
rect -18757 25896 -18725 25930
rect -18824 25840 -18725 25896
rect -4128 25912 -4002 25997
rect -4128 25878 -4069 25912
rect -4035 25878 -4002 25912
rect -4128 25871 -4002 25878
rect -18824 25806 -18791 25840
rect -18757 25806 -18725 25840
rect -18824 25750 -18725 25806
rect -18824 25716 -18791 25750
rect -18757 25716 -18725 25750
rect -18824 25660 -18725 25716
rect -18824 25626 -18791 25660
rect -18757 25626 -18725 25660
rect -18824 25570 -18725 25626
rect -18824 25536 -18791 25570
rect -18757 25536 -18725 25570
rect -18824 25480 -18725 25536
rect -18824 25446 -18791 25480
rect -18757 25446 -18725 25480
rect -18824 25390 -18725 25446
rect -18824 25356 -18791 25390
rect -18757 25356 -18725 25390
rect -18824 25300 -18725 25356
rect -18824 25266 -18791 25300
rect -18757 25266 -18725 25300
rect -18824 25210 -18725 25266
rect -18824 25176 -18791 25210
rect -18757 25176 -18725 25210
rect -18824 25120 -18725 25176
rect -18824 25086 -18791 25120
rect -18757 25086 -18725 25120
rect -18824 25030 -18725 25086
rect -18824 24996 -18791 25030
rect -18757 24996 -18725 25030
rect -18824 24940 -18725 24996
rect -18824 24906 -18791 24940
rect -18757 24906 -18725 24940
rect -18824 24857 -18725 24906
rect -4101 25822 -4002 25871
rect -4101 25788 -4069 25822
rect -4035 25788 -4002 25822
rect -4101 25732 -4002 25788
rect -4101 25698 -4069 25732
rect -4035 25698 -4002 25732
rect -4101 25642 -4002 25698
rect -4101 25608 -4069 25642
rect -4035 25608 -4002 25642
rect -4101 25552 -4002 25608
rect -4101 25518 -4069 25552
rect -4035 25518 -4002 25552
rect -4101 25462 -4002 25518
rect -4101 25428 -4069 25462
rect -4035 25428 -4002 25462
rect -4101 25372 -4002 25428
rect -4101 25338 -4069 25372
rect -4035 25338 -4002 25372
rect -4101 25282 -4002 25338
rect -4101 25248 -4069 25282
rect -4035 25248 -4002 25282
rect -4101 25192 -4002 25248
rect -4101 25158 -4069 25192
rect -4035 25158 -4002 25192
rect -4101 25102 -4002 25158
rect -4101 25068 -4069 25102
rect -4035 25068 -4002 25102
rect -4101 25012 -4002 25068
rect -4101 24978 -4069 25012
rect -4035 24978 -4002 25012
rect -4101 24922 -4002 24978
rect -4101 24888 -4069 24922
rect -4035 24888 -4002 24922
rect -18824 24850 -18698 24857
rect -18824 24816 -18791 24850
rect -18757 24816 -18698 24850
rect -18824 24659 -18698 24816
rect -4101 24832 -4002 24888
rect -4101 24798 -4069 24832
rect -4035 24798 -4002 24832
rect -4101 24781 -4002 24798
rect -18824 24642 -18725 24659
rect -18824 24608 -18791 24642
rect -18757 24608 -18725 24642
rect -18824 24552 -18725 24608
rect -4128 24624 -4002 24781
rect -1712 24718 -1618 30474
rect 4138 24718 4232 30474
rect 29228 28318 29230 28352
rect 30624 28318 30626 28352
rect 32020 28318 32022 28352
rect 33416 28318 33418 28352
rect 34810 28318 34814 28352
rect 36206 28318 36210 28352
rect 37602 28318 37606 28352
rect 38998 28318 39002 28352
rect 40392 28318 40398 28352
rect 41788 28318 41794 28352
rect 43184 28318 43190 28352
rect 44580 28318 44586 28352
rect 45974 28318 45982 28352
rect 47370 28318 47378 28352
rect 48766 28318 48774 28352
rect 50162 28318 50170 28352
rect 29132 27208 29134 28256
rect 30338 27208 30340 28256
rect 30528 27208 30530 28256
rect 31734 27208 31736 28256
rect 31924 27208 31926 28256
rect 33130 27208 33132 28256
rect 33320 27208 33322 28256
rect 34526 27208 34528 28256
rect 34714 27208 34718 28256
rect 35920 27208 35924 28256
rect 36110 27208 36114 28256
rect 37316 27208 37320 28256
rect 37506 27208 37510 28256
rect 38712 27208 38716 28256
rect 38902 27208 38906 28256
rect 40108 27208 40112 28256
rect 40296 27208 40302 28256
rect 41502 27208 41508 28256
rect 41692 27208 41698 28256
rect 42898 27208 42904 28256
rect 43088 27208 43094 28256
rect 44294 27208 44300 28256
rect 44484 27208 44490 28256
rect 45690 27208 45696 28256
rect 45878 27208 45886 28256
rect 47084 27208 47092 28256
rect 47274 27208 47282 28256
rect 48480 27208 48488 28256
rect 48670 27208 48678 28256
rect 49876 27208 49884 28256
rect 50066 27208 50074 28256
rect 51272 27208 51280 28256
rect 29228 27112 29230 27146
rect 30624 27112 30626 27146
rect 32020 27112 32022 27146
rect 33416 27112 33418 27146
rect 34810 27112 34814 27146
rect 36206 27112 36210 27146
rect 37602 27112 37606 27146
rect 38998 27112 39002 27146
rect 40392 27112 40398 27146
rect 41788 27112 41794 27146
rect 43184 27112 43190 27146
rect 44580 27112 44586 27146
rect 45974 27112 45982 27146
rect 47370 27112 47378 27146
rect 48766 27112 48774 27146
rect 50162 27112 50170 27146
rect 29228 26922 29230 26956
rect 30624 26922 30626 26956
rect 32020 26922 32022 26956
rect 33416 26922 33418 26956
rect 34810 26922 34814 26956
rect 36206 26922 36210 26956
rect 37602 26922 37606 26956
rect 38998 26922 39002 26956
rect 40392 26922 40398 26956
rect 41788 26922 41794 26956
rect 43184 26922 43190 26956
rect 44580 26922 44586 26956
rect 45974 26922 45982 26956
rect 47370 26922 47378 26956
rect 48766 26922 48774 26956
rect 50162 26922 50170 26956
rect 29132 25812 29134 26860
rect 30338 25812 30340 26860
rect 30528 25812 30530 26860
rect 31734 25812 31736 26860
rect 31924 25812 31926 26860
rect 33130 25812 33132 26860
rect 33320 25812 33322 26860
rect 34526 25812 34528 26860
rect 34714 25812 34718 26860
rect 35920 25812 35924 26860
rect 36110 25812 36114 26860
rect 37316 25812 37320 26860
rect 37506 25812 37510 26860
rect 38712 25812 38716 26860
rect 38902 25812 38906 26860
rect 40108 25812 40112 26860
rect 40296 25812 40302 26860
rect 41502 25812 41508 26860
rect 41692 25812 41698 26860
rect 42898 25812 42904 26860
rect 43088 25812 43094 26860
rect 44294 25812 44300 26860
rect 44484 25812 44490 26860
rect 45690 25812 45696 26860
rect 45878 25812 45886 26860
rect 47084 25812 47092 26860
rect 47274 25812 47282 26860
rect 48480 25812 48488 26860
rect 48670 25812 48678 26860
rect 49876 25812 49884 26860
rect 50066 25812 50074 26860
rect 51272 25812 51280 26860
rect 29228 25716 29230 25750
rect 30624 25716 30626 25750
rect 32020 25716 32022 25750
rect 33416 25716 33418 25750
rect 34810 25716 34814 25750
rect 36206 25716 36210 25750
rect 37602 25716 37606 25750
rect 38998 25716 39002 25750
rect 40392 25716 40398 25750
rect 41788 25716 41794 25750
rect 43184 25716 43190 25750
rect 44580 25716 44586 25750
rect 45974 25716 45982 25750
rect 47370 25716 47378 25750
rect 48766 25716 48774 25750
rect 50162 25716 50170 25750
rect -1712 24624 4232 24718
rect -4128 24590 -4069 24624
rect -4035 24590 -4002 24624
rect -4128 24583 -4002 24590
rect -18824 24518 -18791 24552
rect -18757 24518 -18725 24552
rect -18824 24462 -18725 24518
rect -18824 24428 -18791 24462
rect -18757 24428 -18725 24462
rect -18824 24372 -18725 24428
rect -18824 24338 -18791 24372
rect -18757 24338 -18725 24372
rect -18824 24282 -18725 24338
rect -18824 24248 -18791 24282
rect -18757 24248 -18725 24282
rect -18824 24192 -18725 24248
rect -18824 24158 -18791 24192
rect -18757 24158 -18725 24192
rect -18824 24102 -18725 24158
rect -18824 24068 -18791 24102
rect -18757 24068 -18725 24102
rect -18824 24012 -18725 24068
rect -18824 23978 -18791 24012
rect -18757 23978 -18725 24012
rect -18824 23922 -18725 23978
rect -18824 23888 -18791 23922
rect -18757 23888 -18725 23922
rect -18824 23832 -18725 23888
rect -18824 23798 -18791 23832
rect -18757 23798 -18725 23832
rect -18824 23742 -18725 23798
rect -18824 23708 -18791 23742
rect -18757 23708 -18725 23742
rect -18824 23652 -18725 23708
rect -18824 23618 -18791 23652
rect -18757 23618 -18725 23652
rect -18824 23569 -18725 23618
rect -4101 24534 -4002 24583
rect -4101 24500 -4069 24534
rect -4035 24500 -4002 24534
rect -4101 24444 -4002 24500
rect -4101 24410 -4069 24444
rect -4035 24410 -4002 24444
rect -4101 24354 -4002 24410
rect -4101 24320 -4069 24354
rect -4035 24320 -4002 24354
rect -4101 24264 -4002 24320
rect -4101 24230 -4069 24264
rect -4035 24230 -4002 24264
rect -4101 24174 -4002 24230
rect -4101 24140 -4069 24174
rect -4035 24140 -4002 24174
rect -4101 24084 -4002 24140
rect -4101 24050 -4069 24084
rect -4035 24050 -4002 24084
rect -4101 23994 -4002 24050
rect 3698 24414 4098 24624
rect 3698 24054 3718 24414
rect 4078 24054 4098 24414
rect 3698 24034 4098 24054
rect -4101 23960 -4069 23994
rect -4035 23960 -4002 23994
rect -4101 23904 -4002 23960
rect -4101 23870 -4069 23904
rect -4035 23870 -4002 23904
rect -4101 23814 -4002 23870
rect -4101 23780 -4069 23814
rect -4035 23780 -4002 23814
rect -4101 23724 -4002 23780
rect -4101 23690 -4069 23724
rect -4035 23690 -4002 23724
rect -4101 23634 -4002 23690
rect -4101 23600 -4069 23634
rect -4035 23600 -4002 23634
rect -18824 23562 -18698 23569
rect -18824 23528 -18791 23562
rect -18757 23528 -18698 23562
rect -18824 23371 -18698 23528
rect -4101 23544 -4002 23600
rect -4101 23510 -4069 23544
rect -4035 23510 -4002 23544
rect -4101 23493 -4002 23510
rect -18824 23354 -18725 23371
rect -18824 23320 -18791 23354
rect -18757 23320 -18725 23354
rect -18824 23264 -18725 23320
rect -4128 23336 -4002 23493
rect -4128 23302 -4069 23336
rect -4035 23302 -4002 23336
rect -4128 23295 -4002 23302
rect -18824 23230 -18791 23264
rect -18757 23230 -18725 23264
rect -18824 23174 -18725 23230
rect -18824 23140 -18791 23174
rect -18757 23140 -18725 23174
rect -18824 23084 -18725 23140
rect -18824 23050 -18791 23084
rect -18757 23050 -18725 23084
rect -18824 22994 -18725 23050
rect -18824 22960 -18791 22994
rect -18757 22960 -18725 22994
rect -18824 22904 -18725 22960
rect -18824 22870 -18791 22904
rect -18757 22870 -18725 22904
rect -18824 22814 -18725 22870
rect -18824 22780 -18791 22814
rect -18757 22780 -18725 22814
rect -18824 22724 -18725 22780
rect -18824 22690 -18791 22724
rect -18757 22690 -18725 22724
rect -18824 22634 -18725 22690
rect -18824 22600 -18791 22634
rect -18757 22600 -18725 22634
rect -18824 22544 -18725 22600
rect -18824 22510 -18791 22544
rect -18757 22510 -18725 22544
rect -18824 22454 -18725 22510
rect -18824 22420 -18791 22454
rect -18757 22420 -18725 22454
rect -18824 22364 -18725 22420
rect -18824 22330 -18791 22364
rect -18757 22330 -18725 22364
rect -18824 22281 -18725 22330
rect -4101 23246 -4002 23295
rect -4101 23212 -4069 23246
rect -4035 23212 -4002 23246
rect -4101 23156 -4002 23212
rect -4101 23122 -4069 23156
rect -4035 23122 -4002 23156
rect -4101 23066 -4002 23122
rect -4101 23032 -4069 23066
rect -4035 23032 -4002 23066
rect -4101 22976 -4002 23032
rect -4101 22942 -4069 22976
rect -4035 22942 -4002 22976
rect -4101 22886 -4002 22942
rect -4101 22852 -4069 22886
rect -4035 22852 -4002 22886
rect -4101 22796 -4002 22852
rect -4101 22762 -4069 22796
rect -4035 22762 -4002 22796
rect -4101 22706 -4002 22762
rect -4101 22672 -4069 22706
rect -4035 22672 -4002 22706
rect -4101 22616 -4002 22672
rect -4101 22582 -4069 22616
rect -4035 22582 -4002 22616
rect -4101 22526 -4002 22582
rect -4101 22492 -4069 22526
rect -4035 22492 -4002 22526
rect -4101 22436 -4002 22492
rect -4101 22402 -4069 22436
rect -4035 22402 -4002 22436
rect -4101 22346 -4002 22402
rect -4101 22312 -4069 22346
rect -4035 22312 -4002 22346
rect -18824 22274 -18698 22281
rect -18824 22240 -18791 22274
rect -18757 22240 -18698 22274
rect -18824 22083 -18698 22240
rect -4101 22256 -4002 22312
rect -4101 22222 -4069 22256
rect -4035 22222 -4002 22256
rect -4101 22205 -4002 22222
rect -18824 22066 -18725 22083
rect -18824 22032 -18791 22066
rect -18757 22032 -18725 22066
rect -18824 21976 -18725 22032
rect -4128 22048 -4002 22205
rect -4128 22014 -4069 22048
rect -4035 22014 -4002 22048
rect -4128 22007 -4002 22014
rect -18824 21942 -18791 21976
rect -18757 21942 -18725 21976
rect -18824 21886 -18725 21942
rect -18824 21852 -18791 21886
rect -18757 21852 -18725 21886
rect -18824 21796 -18725 21852
rect -18824 21762 -18791 21796
rect -18757 21762 -18725 21796
rect -18824 21706 -18725 21762
rect -18824 21672 -18791 21706
rect -18757 21672 -18725 21706
rect -18824 21616 -18725 21672
rect -18824 21582 -18791 21616
rect -18757 21582 -18725 21616
rect -18824 21526 -18725 21582
rect -18824 21492 -18791 21526
rect -18757 21492 -18725 21526
rect -18824 21436 -18725 21492
rect -18824 21402 -18791 21436
rect -18757 21402 -18725 21436
rect -18824 21346 -18725 21402
rect -18824 21312 -18791 21346
rect -18757 21312 -18725 21346
rect -18824 21256 -18725 21312
rect -18824 21222 -18791 21256
rect -18757 21222 -18725 21256
rect -18824 21166 -18725 21222
rect -18824 21132 -18791 21166
rect -18757 21132 -18725 21166
rect -18824 21076 -18725 21132
rect -18824 21042 -18791 21076
rect -18757 21042 -18725 21076
rect -18824 20993 -18725 21042
rect -4101 21958 -4002 22007
rect -4101 21924 -4069 21958
rect -4035 21924 -4002 21958
rect -4101 21868 -4002 21924
rect -4101 21834 -4069 21868
rect -4035 21834 -4002 21868
rect -4101 21778 -4002 21834
rect -4101 21744 -4069 21778
rect -4035 21744 -4002 21778
rect -4101 21688 -4002 21744
rect -4101 21654 -4069 21688
rect -4035 21654 -4002 21688
rect -4101 21598 -4002 21654
rect -4101 21564 -4069 21598
rect -4035 21564 -4002 21598
rect -4101 21508 -4002 21564
rect -4101 21474 -4069 21508
rect -4035 21474 -4002 21508
rect -4101 21418 -4002 21474
rect -4101 21384 -4069 21418
rect -4035 21384 -4002 21418
rect -4101 21328 -4002 21384
rect -4101 21294 -4069 21328
rect -4035 21294 -4002 21328
rect -4101 21238 -4002 21294
rect -4101 21204 -4069 21238
rect -4035 21204 -4002 21238
rect -4101 21148 -4002 21204
rect -4101 21114 -4069 21148
rect -4035 21114 -4002 21148
rect -4101 21058 -4002 21114
rect -4101 21024 -4069 21058
rect -4035 21024 -4002 21058
rect -18824 20986 -18698 20993
rect -18824 20952 -18791 20986
rect -18757 20952 -18698 20986
rect -18824 20795 -18698 20952
rect -4101 20968 -4002 21024
rect -4101 20934 -4069 20968
rect -4035 20934 -4002 20968
rect -4101 20917 -4002 20934
rect -18824 20778 -18725 20795
rect -18824 20744 -18791 20778
rect -18757 20744 -18725 20778
rect -18824 20688 -18725 20744
rect -4128 20760 -4002 20917
rect -4128 20726 -4069 20760
rect -4035 20726 -4002 20760
rect -4128 20719 -4002 20726
rect -18824 20654 -18791 20688
rect -18757 20654 -18725 20688
rect -18824 20598 -18725 20654
rect -18824 20564 -18791 20598
rect -18757 20564 -18725 20598
rect -18824 20508 -18725 20564
rect -18824 20474 -18791 20508
rect -18757 20474 -18725 20508
rect -18824 20418 -18725 20474
rect -18824 20384 -18791 20418
rect -18757 20384 -18725 20418
rect -18824 20328 -18725 20384
rect -18824 20294 -18791 20328
rect -18757 20294 -18725 20328
rect -18824 20238 -18725 20294
rect -18824 20204 -18791 20238
rect -18757 20204 -18725 20238
rect -18824 20148 -18725 20204
rect -18824 20114 -18791 20148
rect -18757 20114 -18725 20148
rect -18824 20058 -18725 20114
rect -18824 20024 -18791 20058
rect -18757 20024 -18725 20058
rect -18824 19968 -18725 20024
rect -18824 19934 -18791 19968
rect -18757 19934 -18725 19968
rect -18824 19878 -18725 19934
rect -18824 19844 -18791 19878
rect -18757 19844 -18725 19878
rect -18824 19788 -18725 19844
rect -18824 19754 -18791 19788
rect -18757 19754 -18725 19788
rect -18824 19705 -18725 19754
rect -4101 20670 -4002 20719
rect -4101 20636 -4069 20670
rect -4035 20636 -4002 20670
rect -4101 20580 -4002 20636
rect -4101 20546 -4069 20580
rect -4035 20546 -4002 20580
rect -4101 20490 -4002 20546
rect -4101 20456 -4069 20490
rect -4035 20456 -4002 20490
rect -4101 20400 -4002 20456
rect -4101 20366 -4069 20400
rect -4035 20366 -4002 20400
rect -4101 20310 -4002 20366
rect -4101 20276 -4069 20310
rect -4035 20276 -4002 20310
rect -4101 20220 -4002 20276
rect -4101 20186 -4069 20220
rect -4035 20186 -4002 20220
rect -4101 20130 -4002 20186
rect -4101 20096 -4069 20130
rect -4035 20096 -4002 20130
rect -4101 20040 -4002 20096
rect -4101 20006 -4069 20040
rect -4035 20006 -4002 20040
rect -4101 19950 -4002 20006
rect -4101 19916 -4069 19950
rect -4035 19916 -4002 19950
rect -4101 19860 -4002 19916
rect -4101 19826 -4069 19860
rect -4035 19826 -4002 19860
rect -4101 19770 -4002 19826
rect -4101 19736 -4069 19770
rect -4035 19736 -4002 19770
rect -18824 19698 -18698 19705
rect -18824 19664 -18791 19698
rect -18757 19664 -18698 19698
rect -18824 19507 -18698 19664
rect -4101 19680 -4002 19736
rect -4101 19646 -4069 19680
rect -4035 19646 -4002 19680
rect -4101 19629 -4002 19646
rect -18824 19490 -18725 19507
rect -18824 19456 -18791 19490
rect -18757 19456 -18725 19490
rect -18824 19400 -18725 19456
rect -4128 19472 -4002 19629
rect -4128 19438 -4069 19472
rect -4035 19438 -4002 19472
rect -4128 19431 -4002 19438
rect -18824 19366 -18791 19400
rect -18757 19366 -18725 19400
rect -18824 19310 -18725 19366
rect -18824 19276 -18791 19310
rect -18757 19276 -18725 19310
rect -18824 19220 -18725 19276
rect -18824 19186 -18791 19220
rect -18757 19186 -18725 19220
rect -18824 19130 -18725 19186
rect -18824 19096 -18791 19130
rect -18757 19096 -18725 19130
rect -18824 19040 -18725 19096
rect -18824 19006 -18791 19040
rect -18757 19006 -18725 19040
rect -18824 18950 -18725 19006
rect -18824 18916 -18791 18950
rect -18757 18916 -18725 18950
rect -18824 18860 -18725 18916
rect -18824 18826 -18791 18860
rect -18757 18826 -18725 18860
rect -18824 18770 -18725 18826
rect -18824 18736 -18791 18770
rect -18757 18736 -18725 18770
rect -18824 18680 -18725 18736
rect -18824 18646 -18791 18680
rect -18757 18646 -18725 18680
rect -18824 18590 -18725 18646
rect -18824 18556 -18791 18590
rect -18757 18556 -18725 18590
rect -18824 18500 -18725 18556
rect -18824 18466 -18791 18500
rect -18757 18466 -18725 18500
rect -18824 18417 -18725 18466
rect -4101 19382 -4002 19431
rect -4101 19348 -4069 19382
rect -4035 19348 -4002 19382
rect -4101 19292 -4002 19348
rect -4101 19258 -4069 19292
rect -4035 19258 -4002 19292
rect -4101 19202 -4002 19258
rect -4101 19168 -4069 19202
rect -4035 19168 -4002 19202
rect -4101 19112 -4002 19168
rect -4101 19078 -4069 19112
rect -4035 19078 -4002 19112
rect -4101 19048 -4002 19078
rect -4101 19022 -2560 19048
rect -4101 18988 -4069 19022
rect -4035 19016 -2560 19022
rect -4035 18988 -2944 19016
rect -4101 18932 -2944 18988
rect -4101 18898 -4069 18932
rect -4035 18898 -2944 18932
rect -4101 18842 -2944 18898
rect -4101 18808 -4069 18842
rect -4035 18808 -2944 18842
rect -4101 18752 -2944 18808
rect -4101 18718 -4069 18752
rect -4035 18718 -2944 18752
rect -4101 18664 -2944 18718
rect -2592 18664 -2560 19016
rect -4101 18662 -2560 18664
rect -4101 18628 -4069 18662
rect -4035 18630 -2560 18662
rect -4035 18628 -4002 18630
rect -4101 18572 -4002 18628
rect -4101 18538 -4069 18572
rect -4035 18538 -4002 18572
rect -4101 18482 -4002 18538
rect -4101 18448 -4069 18482
rect -4035 18448 -4002 18482
rect -18824 18410 -18698 18417
rect -18824 18376 -18791 18410
rect -18757 18376 -18698 18410
rect -18824 18219 -18698 18376
rect -4101 18392 -4002 18448
rect -4101 18358 -4069 18392
rect -4035 18358 -4002 18392
rect -4101 18341 -4002 18358
rect -18824 18202 -18725 18219
rect -18824 18168 -18791 18202
rect -18757 18168 -18725 18202
rect -18824 18112 -18725 18168
rect -4128 18184 -4002 18341
rect -4128 18150 -4069 18184
rect -4035 18150 -4002 18184
rect -4128 18143 -4002 18150
rect -18824 18078 -18791 18112
rect -18757 18078 -18725 18112
rect -18824 18022 -18725 18078
rect -18824 17988 -18791 18022
rect -18757 17988 -18725 18022
rect -18824 17932 -18725 17988
rect -18824 17898 -18791 17932
rect -18757 17898 -18725 17932
rect -18824 17842 -18725 17898
rect -18824 17808 -18791 17842
rect -18757 17808 -18725 17842
rect -18824 17752 -18725 17808
rect -18824 17718 -18791 17752
rect -18757 17718 -18725 17752
rect -18824 17662 -18725 17718
rect -18824 17628 -18791 17662
rect -18757 17628 -18725 17662
rect -18824 17572 -18725 17628
rect -18824 17538 -18791 17572
rect -18757 17538 -18725 17572
rect -18824 17482 -18725 17538
rect -18824 17448 -18791 17482
rect -18757 17448 -18725 17482
rect -18824 17392 -18725 17448
rect -18824 17358 -18791 17392
rect -18757 17358 -18725 17392
rect -18824 17302 -18725 17358
rect -18824 17268 -18791 17302
rect -18757 17268 -18725 17302
rect -18824 17212 -18725 17268
rect -18824 17178 -18791 17212
rect -18757 17178 -18725 17212
rect -18824 17129 -18725 17178
rect -4101 18094 -4002 18143
rect -4101 18060 -4069 18094
rect -4035 18060 -4002 18094
rect -4101 18004 -4002 18060
rect -4101 17970 -4069 18004
rect -4035 17970 -4002 18004
rect -4101 17914 -4002 17970
rect -4101 17880 -4069 17914
rect -4035 17880 -4002 17914
rect -4101 17824 -4002 17880
rect -4101 17790 -4069 17824
rect -4035 17790 -4002 17824
rect -4101 17734 -4002 17790
rect -4101 17700 -4069 17734
rect -4035 17700 -4002 17734
rect -4101 17644 -4002 17700
rect -4101 17610 -4069 17644
rect -4035 17610 -4002 17644
rect -4101 17554 -4002 17610
rect -4101 17520 -4069 17554
rect -4035 17520 -4002 17554
rect -4101 17464 -4002 17520
rect -4101 17430 -4069 17464
rect -4035 17430 -4002 17464
rect -4101 17374 -4002 17430
rect -4101 17340 -4069 17374
rect -4035 17340 -4002 17374
rect -4101 17284 -4002 17340
rect -4101 17250 -4069 17284
rect -4035 17250 -4002 17284
rect -4101 17194 -4002 17250
rect -4101 17160 -4069 17194
rect -4035 17160 -4002 17194
rect -18824 17122 -18698 17129
rect -18824 17088 -18791 17122
rect -18757 17088 -18698 17122
rect -18824 17003 -18698 17088
rect -4101 17104 -4002 17160
rect -4101 17070 -4069 17104
rect -4035 17070 -4002 17104
rect -4101 17053 -4002 17070
rect -18824 16986 -18725 17003
rect -18824 16952 -18791 16986
rect -18757 16952 -18725 16986
rect -18824 16896 -18725 16952
rect -18824 16862 -18791 16896
rect -18757 16862 -18725 16896
rect -18824 16806 -18725 16862
rect -4128 16896 -4002 17053
rect -4128 16862 -4069 16896
rect -4035 16862 -4002 16896
rect -4128 16855 -4002 16862
rect -18824 16772 -18791 16806
rect -18757 16772 -18725 16806
rect -18824 16716 -18725 16772
rect -18824 16682 -18791 16716
rect -18757 16682 -18725 16716
rect -18824 16626 -18725 16682
rect -18824 16592 -18791 16626
rect -18757 16592 -18725 16626
rect -18824 16536 -18725 16592
rect -18824 16502 -18791 16536
rect -18757 16502 -18725 16536
rect -18824 16446 -18725 16502
rect -18824 16412 -18791 16446
rect -18757 16412 -18725 16446
rect -18824 16356 -18725 16412
rect -18824 16322 -18791 16356
rect -18757 16322 -18725 16356
rect -18824 16266 -18725 16322
rect -18824 16232 -18791 16266
rect -18757 16232 -18725 16266
rect -18824 16176 -18725 16232
rect -18824 16142 -18791 16176
rect -18757 16142 -18725 16176
rect -18824 16086 -18725 16142
rect -18824 16052 -18791 16086
rect -18757 16052 -18725 16086
rect -18824 15996 -18725 16052
rect -18824 15962 -18791 15996
rect -18757 15962 -18725 15996
rect -18824 15913 -18725 15962
rect -4101 16806 -4002 16855
rect -4101 16772 -4069 16806
rect -4035 16772 -4002 16806
rect -4101 16716 -4002 16772
rect -4101 16682 -4069 16716
rect -4035 16682 -4002 16716
rect -4101 16626 -4002 16682
rect -4101 16592 -4069 16626
rect -4035 16592 -4002 16626
rect -4101 16536 -4002 16592
rect -4101 16502 -4069 16536
rect -4035 16502 -4002 16536
rect -4101 16446 -4002 16502
rect -4101 16412 -4069 16446
rect -4035 16412 -4002 16446
rect -4101 16356 -4002 16412
rect -4101 16322 -4069 16356
rect -4035 16322 -4002 16356
rect -4101 16266 -4002 16322
rect -4101 16232 -4069 16266
rect -4035 16232 -4002 16266
rect -4101 16176 -4002 16232
rect -4101 16142 -4069 16176
rect -4035 16142 -4002 16176
rect -4101 16086 -4002 16142
rect -4101 16052 -4069 16086
rect -4035 16052 -4002 16086
rect -4101 15996 -4002 16052
rect -4101 15962 -4069 15996
rect -4035 15962 -4002 15996
rect -18824 15906 -18698 15913
rect -18824 15872 -18791 15906
rect -18757 15872 -18698 15906
rect -18824 15715 -18698 15872
rect -4101 15906 -4002 15962
rect -4101 15872 -4069 15906
rect -4035 15872 -4002 15906
rect -4101 15816 -4002 15872
rect -4101 15782 -4069 15816
rect -4035 15782 -4002 15816
rect -4101 15765 -4002 15782
rect -18824 15698 -18725 15715
rect -18824 15664 -18791 15698
rect -18757 15664 -18725 15698
rect -18824 15608 -18725 15664
rect -18824 15574 -18791 15608
rect -18757 15574 -18725 15608
rect -18824 15518 -18725 15574
rect -4128 15608 -4002 15765
rect -4128 15574 -4069 15608
rect -4035 15574 -4002 15608
rect -4128 15567 -4002 15574
rect -18824 15484 -18791 15518
rect -18757 15484 -18725 15518
rect -18824 15428 -18725 15484
rect -18824 15394 -18791 15428
rect -18757 15394 -18725 15428
rect -18824 15338 -18725 15394
rect -18824 15304 -18791 15338
rect -18757 15304 -18725 15338
rect -18824 15248 -18725 15304
rect -18824 15214 -18791 15248
rect -18757 15214 -18725 15248
rect -18824 15158 -18725 15214
rect -18824 15124 -18791 15158
rect -18757 15124 -18725 15158
rect -18824 15068 -18725 15124
rect -18824 15034 -18791 15068
rect -18757 15034 -18725 15068
rect -18824 14978 -18725 15034
rect -18824 14944 -18791 14978
rect -18757 14944 -18725 14978
rect -18824 14888 -18725 14944
rect -18824 14854 -18791 14888
rect -18757 14854 -18725 14888
rect -18824 14798 -18725 14854
rect -18824 14764 -18791 14798
rect -18757 14764 -18725 14798
rect -18824 14708 -18725 14764
rect -18824 14674 -18791 14708
rect -18757 14674 -18725 14708
rect -18824 14625 -18725 14674
rect -4101 15518 -4002 15567
rect -4101 15484 -4069 15518
rect -4035 15484 -4002 15518
rect -4101 15428 -4002 15484
rect -4101 15394 -4069 15428
rect -4035 15394 -4002 15428
rect -4101 15338 -4002 15394
rect -4101 15304 -4069 15338
rect -4035 15304 -4002 15338
rect -4101 15248 -4002 15304
rect -4101 15214 -4069 15248
rect -4035 15214 -4002 15248
rect -4101 15158 -4002 15214
rect -4101 15124 -4069 15158
rect -4035 15124 -4002 15158
rect -4101 15068 -4002 15124
rect -4101 15034 -4069 15068
rect -4035 15034 -4002 15068
rect -4101 14978 -4002 15034
rect -4101 14944 -4069 14978
rect -4035 14944 -4002 14978
rect -4101 14888 -4002 14944
rect -4101 14854 -4069 14888
rect -4035 14854 -4002 14888
rect -4101 14798 -4002 14854
rect -4101 14764 -4069 14798
rect -4035 14764 -4002 14798
rect -4101 14708 -4002 14764
rect -4101 14674 -4069 14708
rect -4035 14674 -4002 14708
rect -18824 14618 -18698 14625
rect -18824 14584 -18791 14618
rect -18757 14584 -18698 14618
rect -18824 14427 -18698 14584
rect -4101 14618 -4002 14674
rect -4101 14584 -4069 14618
rect -4035 14584 -4002 14618
rect -4101 14528 -4002 14584
rect -4101 14494 -4069 14528
rect -4035 14494 -4002 14528
rect -4101 14477 -4002 14494
rect -18824 14410 -18725 14427
rect -18824 14376 -18791 14410
rect -18757 14376 -18725 14410
rect -18824 14320 -18725 14376
rect -18824 14286 -18791 14320
rect -18757 14286 -18725 14320
rect -18824 14230 -18725 14286
rect -4128 14320 -4002 14477
rect -4128 14286 -4069 14320
rect -4035 14286 -4002 14320
rect -4128 14279 -4002 14286
rect -18824 14196 -18791 14230
rect -18757 14196 -18725 14230
rect -18824 14140 -18725 14196
rect -18824 14106 -18791 14140
rect -18757 14106 -18725 14140
rect -18824 14050 -18725 14106
rect -18824 14016 -18791 14050
rect -18757 14016 -18725 14050
rect -18824 13960 -18725 14016
rect -18824 13926 -18791 13960
rect -18757 13926 -18725 13960
rect -18824 13870 -18725 13926
rect -18824 13836 -18791 13870
rect -18757 13836 -18725 13870
rect -18824 13780 -18725 13836
rect -18824 13746 -18791 13780
rect -18757 13746 -18725 13780
rect -18824 13690 -18725 13746
rect -18824 13656 -18791 13690
rect -18757 13656 -18725 13690
rect -18824 13600 -18725 13656
rect -18824 13566 -18791 13600
rect -18757 13566 -18725 13600
rect -18824 13510 -18725 13566
rect -18824 13476 -18791 13510
rect -18757 13476 -18725 13510
rect -18824 13420 -18725 13476
rect -18824 13386 -18791 13420
rect -18757 13386 -18725 13420
rect -18824 13337 -18725 13386
rect -4101 14230 -4002 14279
rect -4101 14196 -4069 14230
rect -4035 14196 -4002 14230
rect -4101 14140 -4002 14196
rect -4101 14106 -4069 14140
rect -4035 14106 -4002 14140
rect -4101 14050 -4002 14106
rect -4101 14016 -4069 14050
rect -4035 14016 -4002 14050
rect -4101 13960 -4002 14016
rect -4101 13926 -4069 13960
rect -4035 13926 -4002 13960
rect -4101 13870 -4002 13926
rect -4101 13836 -4069 13870
rect -4035 13836 -4002 13870
rect -4101 13780 -4002 13836
rect -4101 13746 -4069 13780
rect -4035 13746 -4002 13780
rect -4101 13690 -4002 13746
rect -4101 13656 -4069 13690
rect -4035 13656 -4002 13690
rect -4101 13600 -4002 13656
rect -4101 13566 -4069 13600
rect -4035 13566 -4002 13600
rect -4101 13510 -4002 13566
rect -4101 13476 -4069 13510
rect -4035 13476 -4002 13510
rect -4101 13420 -4002 13476
rect -4101 13386 -4069 13420
rect -4035 13386 -4002 13420
rect -18824 13330 -18698 13337
rect -18824 13296 -18791 13330
rect -18757 13296 -18698 13330
rect -18824 13189 -18698 13296
rect -4101 13330 -4002 13386
rect -4101 13296 -4069 13330
rect -4035 13296 -4002 13330
rect -4101 13240 -4002 13296
rect -4101 13216 -4070 13240
rect -18255 13189 -18057 13216
rect -16967 13189 -16769 13216
rect -15679 13189 -15481 13216
rect -14391 13189 -14193 13216
rect -13103 13189 -12905 13216
rect -11815 13189 -11617 13216
rect -10527 13189 -10329 13216
rect -9239 13189 -9041 13216
rect -7951 13189 -7825 13216
rect -6735 13189 -6537 13216
rect -5447 13189 -5249 13216
rect -4104 13206 -4070 13216
rect -4034 13206 -4002 13240
rect -4104 13192 -4002 13206
rect -4159 13189 -4002 13192
rect -18824 13157 -4002 13189
rect -18824 13123 -18788 13157
rect -18754 13123 -18698 13157
rect -18664 13123 -18608 13157
rect -18574 13123 -18518 13157
rect -18484 13123 -18428 13157
rect -18394 13123 -18338 13157
rect -18304 13123 -18248 13157
rect -18214 13123 -18040 13157
rect -18006 13123 -17950 13157
rect -17916 13123 -17860 13157
rect -17826 13123 -17770 13157
rect -17736 13123 -17680 13157
rect -17646 13123 -17590 13157
rect -17556 13123 -17500 13157
rect -17466 13123 -17410 13157
rect -17376 13123 -17320 13157
rect -17286 13123 -17230 13157
rect -17196 13123 -17140 13157
rect -17106 13123 -17050 13157
rect -17016 13123 -16960 13157
rect -16926 13123 -16752 13157
rect -16718 13123 -16662 13157
rect -16628 13123 -16572 13157
rect -16538 13123 -16482 13157
rect -16448 13123 -16392 13157
rect -16358 13123 -16302 13157
rect -16268 13123 -16212 13157
rect -16178 13123 -16122 13157
rect -16088 13123 -16032 13157
rect -15998 13123 -15942 13157
rect -15908 13123 -15852 13157
rect -15818 13123 -15762 13157
rect -15728 13123 -15672 13157
rect -15638 13123 -15464 13157
rect -15430 13123 -15374 13157
rect -15340 13123 -15284 13157
rect -15250 13123 -15194 13157
rect -15160 13123 -15104 13157
rect -15070 13123 -15014 13157
rect -14980 13123 -14924 13157
rect -14890 13123 -14834 13157
rect -14800 13123 -14744 13157
rect -14710 13123 -14654 13157
rect -14620 13123 -14564 13157
rect -14530 13123 -14474 13157
rect -14440 13123 -14384 13157
rect -14350 13123 -14176 13157
rect -14142 13123 -14086 13157
rect -14052 13123 -13996 13157
rect -13962 13123 -13906 13157
rect -13872 13123 -13816 13157
rect -13782 13123 -13726 13157
rect -13692 13123 -13636 13157
rect -13602 13123 -13546 13157
rect -13512 13123 -13456 13157
rect -13422 13123 -13366 13157
rect -13332 13123 -13276 13157
rect -13242 13123 -13186 13157
rect -13152 13123 -13096 13157
rect -13062 13123 -12888 13157
rect -12854 13123 -12798 13157
rect -12764 13123 -12708 13157
rect -12674 13123 -12618 13157
rect -12584 13123 -12528 13157
rect -12494 13123 -12438 13157
rect -12404 13123 -12348 13157
rect -12314 13123 -12258 13157
rect -12224 13123 -12168 13157
rect -12134 13123 -12078 13157
rect -12044 13123 -11988 13157
rect -11954 13123 -11898 13157
rect -11864 13123 -11808 13157
rect -11774 13123 -11600 13157
rect -11566 13123 -11510 13157
rect -11476 13123 -11420 13157
rect -11386 13123 -11330 13157
rect -11296 13123 -11240 13157
rect -11206 13123 -11150 13157
rect -11116 13123 -11060 13157
rect -11026 13123 -10970 13157
rect -10936 13123 -10880 13157
rect -10846 13123 -10790 13157
rect -10756 13123 -10700 13157
rect -10666 13123 -10610 13157
rect -10576 13123 -10520 13157
rect -10486 13123 -10312 13157
rect -10278 13123 -10222 13157
rect -10188 13123 -10132 13157
rect -10098 13123 -10042 13157
rect -10008 13123 -9952 13157
rect -9918 13123 -9862 13157
rect -9828 13123 -9772 13157
rect -9738 13123 -9682 13157
rect -9648 13123 -9592 13157
rect -9558 13123 -9502 13157
rect -9468 13123 -9412 13157
rect -9378 13123 -9322 13157
rect -9288 13123 -9232 13157
rect -9198 13123 -9024 13157
rect -8990 13123 -8934 13157
rect -8900 13123 -8844 13157
rect -8810 13123 -8754 13157
rect -8720 13123 -8664 13157
rect -8630 13123 -8574 13157
rect -8540 13123 -8484 13157
rect -8450 13123 -8394 13157
rect -8360 13123 -8304 13157
rect -8270 13123 -8214 13157
rect -8180 13123 -8124 13157
rect -8090 13123 -8034 13157
rect -8000 13123 -7944 13157
rect -7910 13123 -7808 13157
rect -7774 13123 -7718 13157
rect -7684 13123 -7628 13157
rect -7594 13123 -7538 13157
rect -7504 13123 -7448 13157
rect -7414 13123 -7358 13157
rect -7324 13123 -7268 13157
rect -7234 13123 -7178 13157
rect -7144 13123 -7088 13157
rect -7054 13123 -6998 13157
rect -6964 13123 -6908 13157
rect -6874 13123 -6818 13157
rect -6784 13123 -6728 13157
rect -6694 13123 -6520 13157
rect -6486 13123 -6430 13157
rect -6396 13123 -6340 13157
rect -6306 13123 -6250 13157
rect -6216 13123 -6160 13157
rect -6126 13123 -6070 13157
rect -6036 13123 -5980 13157
rect -5946 13123 -5890 13157
rect -5856 13123 -5800 13157
rect -5766 13123 -5710 13157
rect -5676 13123 -5620 13157
rect -5586 13123 -5530 13157
rect -5496 13123 -5440 13157
rect -5406 13123 -5232 13157
rect -5198 13123 -5142 13157
rect -5108 13123 -5052 13157
rect -5018 13123 -4962 13157
rect -4928 13123 -4872 13157
rect -4838 13123 -4782 13157
rect -4748 13123 -4692 13157
rect -4658 13123 -4602 13157
rect -4568 13123 -4512 13157
rect -4478 13123 -4422 13157
rect -4388 13123 -4332 13157
rect -4298 13123 -4242 13157
rect -4208 13123 -4152 13157
rect -4118 13123 -4002 13157
rect -18824 13090 -4002 13123
rect -18824 13084 -18766 13090
<< viali >>
rect -1358 30276 -310 30310
rect 38 30276 1086 30310
rect 1434 30276 2482 30310
rect 2830 30276 3878 30310
rect -1454 29166 -1420 30214
rect -248 29166 -214 30214
rect -58 29166 -24 30214
rect 1148 29166 1182 30214
rect 1338 29166 1372 30214
rect 2544 29166 2578 30214
rect 2734 29166 2768 30214
rect 3940 29166 3974 30214
rect -1358 29070 -310 29104
rect 38 29070 1086 29104
rect 1434 29070 2482 29104
rect 2830 29070 3878 29104
rect -1358 28880 -310 28914
rect 38 28880 1086 28914
rect 1434 28880 2482 28914
rect 2830 28880 3878 28914
rect -1454 27770 -1420 28818
rect -248 27770 -214 28818
rect -58 27770 -24 28818
rect 1148 27770 1182 28818
rect 1338 27770 1372 28818
rect 2544 27770 2578 28818
rect 2734 27770 2768 28818
rect 3940 27770 3974 28818
rect -1358 27674 -310 27708
rect 38 27674 1086 27708
rect 1434 27674 2482 27708
rect 2830 27674 3878 27708
rect -1358 27484 -310 27518
rect 38 27484 1086 27518
rect 1434 27484 2482 27518
rect 2830 27484 3878 27518
rect -1454 26374 -1420 27422
rect -248 26374 -214 27422
rect -58 26374 -24 27422
rect 1148 26374 1182 27422
rect 1338 26374 1372 27422
rect 2544 26374 2578 27422
rect 2734 26374 2768 27422
rect 3940 26374 3974 27422
rect -1358 26278 -310 26312
rect 38 26278 1086 26312
rect 1434 26278 2482 26312
rect 2830 26278 3878 26312
rect -1358 26088 -310 26122
rect 38 26088 1086 26122
rect 1434 26088 2482 26122
rect 2830 26088 3878 26122
rect -1454 24978 -1420 26026
rect -248 24978 -214 26026
rect -58 24978 -24 26026
rect 1148 24978 1182 26026
rect 1338 24978 1372 26026
rect 2544 24978 2578 26026
rect 2734 24978 2768 26026
rect 3940 24978 3974 26026
rect -1358 24882 -310 24916
rect 38 24882 1086 24916
rect 1434 24882 2482 24916
rect 2830 24882 3878 24916
rect 9476 28528 51428 28562
rect 9380 25602 9414 28466
rect 9686 28318 10734 28352
rect 11082 28318 12130 28352
rect 12478 28318 13526 28352
rect 13874 28318 14922 28352
rect 15270 28318 16318 28352
rect 16666 28318 17714 28352
rect 18062 28318 19110 28352
rect 19458 28318 20506 28352
rect 20854 28318 21902 28352
rect 22250 28318 23298 28352
rect 23646 28318 24694 28352
rect 25042 28318 26090 28352
rect 26438 28318 27486 28352
rect 27834 28318 28882 28352
rect 29230 28318 30278 28352
rect 30626 28318 31674 28352
rect 32022 28318 33070 28352
rect 33418 28318 34466 28352
rect 34814 28318 35862 28352
rect 36210 28318 37258 28352
rect 37606 28318 38654 28352
rect 39002 28318 40050 28352
rect 40398 28318 41446 28352
rect 41794 28318 42842 28352
rect 43190 28318 44238 28352
rect 44586 28318 45634 28352
rect 45982 28318 47030 28352
rect 47378 28318 48426 28352
rect 48774 28318 49822 28352
rect 50170 28318 51218 28352
rect 9590 27208 9624 28256
rect 10796 27208 10830 28256
rect 10986 27208 11020 28256
rect 12192 27208 12226 28256
rect 12382 27208 12416 28256
rect 13588 27208 13622 28256
rect 13778 27208 13812 28256
rect 14984 27208 15018 28256
rect 15174 27208 15208 28256
rect 16380 27208 16414 28256
rect 16570 27208 16604 28256
rect 17776 27208 17810 28256
rect 17966 27208 18000 28256
rect 19172 27208 19206 28256
rect 19362 27208 19396 28256
rect 20568 27208 20602 28256
rect 20758 27208 20792 28256
rect 21964 27208 21998 28256
rect 22154 27208 22188 28256
rect 23360 27208 23394 28256
rect 23550 27208 23584 28256
rect 24756 27208 24790 28256
rect 24946 27208 24980 28256
rect 26152 27208 26186 28256
rect 26342 27208 26376 28256
rect 27548 27208 27582 28256
rect 27738 27208 27772 28256
rect 28944 27208 28978 28256
rect 29134 27208 29168 28256
rect 30340 27208 30374 28256
rect 30530 27208 30564 28256
rect 31736 27208 31770 28256
rect 31926 27208 31960 28256
rect 33132 27208 33166 28256
rect 33322 27208 33356 28256
rect 34528 27208 34562 28256
rect 34718 27208 34752 28256
rect 35924 27208 35958 28256
rect 36114 27208 36148 28256
rect 37320 27208 37354 28256
rect 37510 27208 37544 28256
rect 38716 27208 38750 28256
rect 38906 27208 38940 28256
rect 40112 27208 40146 28256
rect 40302 27208 40336 28256
rect 41508 27208 41542 28256
rect 41698 27208 41732 28256
rect 42904 27208 42938 28256
rect 43094 27208 43128 28256
rect 44300 27208 44334 28256
rect 44490 27208 44524 28256
rect 45696 27208 45730 28256
rect 45886 27208 45920 28256
rect 47092 27208 47126 28256
rect 47282 27208 47316 28256
rect 48488 27208 48522 28256
rect 48678 27208 48712 28256
rect 49884 27208 49918 28256
rect 50074 27208 50108 28256
rect 51280 27208 51314 28256
rect 9686 27112 9786 27146
rect 10634 27112 10734 27146
rect 11082 27112 11182 27146
rect 12030 27112 12130 27146
rect 12478 27112 12578 27146
rect 13426 27112 13526 27146
rect 13874 27112 13974 27146
rect 14822 27112 14922 27146
rect 15270 27112 15370 27146
rect 16218 27112 16318 27146
rect 16666 27112 16766 27146
rect 17614 27112 17714 27146
rect 18062 27112 18162 27146
rect 19010 27112 19110 27146
rect 19458 27112 19558 27146
rect 20406 27112 20506 27146
rect 20854 27112 20954 27146
rect 21802 27112 21902 27146
rect 22250 27112 22350 27146
rect 23198 27112 23298 27146
rect 23646 27112 23746 27146
rect 24594 27112 24694 27146
rect 25042 27112 25142 27146
rect 25990 27112 26090 27146
rect 26438 27112 26538 27146
rect 27386 27112 27486 27146
rect 27834 27112 27934 27146
rect 28782 27112 28882 27146
rect 29230 27112 29330 27146
rect 30178 27112 30278 27146
rect 30626 27112 30726 27146
rect 31574 27112 31674 27146
rect 32022 27112 32122 27146
rect 32970 27112 33070 27146
rect 33418 27112 33518 27146
rect 34366 27112 34466 27146
rect 34814 27112 34914 27146
rect 35762 27112 35862 27146
rect 36210 27112 36310 27146
rect 37158 27112 37258 27146
rect 37606 27112 37706 27146
rect 38554 27112 38654 27146
rect 39002 27112 39102 27146
rect 39950 27112 40050 27146
rect 40398 27112 40498 27146
rect 41346 27112 41446 27146
rect 41794 27112 41894 27146
rect 42742 27112 42842 27146
rect 43190 27112 43290 27146
rect 44138 27112 44238 27146
rect 44586 27112 44686 27146
rect 45534 27112 45634 27146
rect 45982 27112 46082 27146
rect 46930 27112 47030 27146
rect 47378 27112 47478 27146
rect 48326 27112 48426 27146
rect 48774 27112 48874 27146
rect 49722 27112 49822 27146
rect 50170 27112 50270 27146
rect 51118 27112 51218 27146
rect 9686 26922 9786 26956
rect 10634 26922 10734 26956
rect 11082 26922 11182 26956
rect 12030 26922 12130 26956
rect 12478 26922 12578 26956
rect 13426 26922 13526 26956
rect 13874 26922 13974 26956
rect 14822 26922 14922 26956
rect 15270 26922 15370 26956
rect 16218 26922 16318 26956
rect 16666 26922 16766 26956
rect 17614 26922 17714 26956
rect 18062 26922 18162 26956
rect 19010 26922 19110 26956
rect 19458 26922 19558 26956
rect 20406 26922 20506 26956
rect 20854 26922 20954 26956
rect 21802 26922 21902 26956
rect 22250 26922 22350 26956
rect 23198 26922 23298 26956
rect 23646 26922 23746 26956
rect 24594 26922 24694 26956
rect 25042 26922 25142 26956
rect 25990 26922 26090 26956
rect 26438 26922 26538 26956
rect 27386 26922 27486 26956
rect 27834 26922 27934 26956
rect 28782 26922 28882 26956
rect 29230 26922 29330 26956
rect 30178 26922 30278 26956
rect 30626 26922 30726 26956
rect 31574 26922 31674 26956
rect 32022 26922 32122 26956
rect 32970 26922 33070 26956
rect 33418 26922 33518 26956
rect 34366 26922 34466 26956
rect 34814 26922 34914 26956
rect 35762 26922 35862 26956
rect 36210 26922 36310 26956
rect 37158 26922 37258 26956
rect 37606 26922 37706 26956
rect 38554 26922 38654 26956
rect 39002 26922 39102 26956
rect 39950 26922 40050 26956
rect 40398 26922 40498 26956
rect 41346 26922 41446 26956
rect 41794 26922 41894 26956
rect 42742 26922 42842 26956
rect 43190 26922 43290 26956
rect 44138 26922 44238 26956
rect 44586 26922 44686 26956
rect 45534 26922 45634 26956
rect 45982 26922 46082 26956
rect 46930 26922 47030 26956
rect 47378 26922 47478 26956
rect 48326 26922 48426 26956
rect 48774 26922 48874 26956
rect 49722 26922 49822 26956
rect 50170 26922 50270 26956
rect 51118 26922 51218 26956
rect 9590 25812 9624 26860
rect 10796 25812 10830 26860
rect 10986 25812 11020 26860
rect 12192 25812 12226 26860
rect 12382 25812 12416 26860
rect 13588 25812 13622 26860
rect 13778 25812 13812 26860
rect 14984 25812 15018 26860
rect 15174 25812 15208 26860
rect 16380 25812 16414 26860
rect 16570 25812 16604 26860
rect 17776 25812 17810 26860
rect 17966 25812 18000 26860
rect 19172 25812 19206 26860
rect 19362 25812 19396 26860
rect 20568 25812 20602 26860
rect 20758 25812 20792 26860
rect 21964 25812 21998 26860
rect 22154 25812 22188 26860
rect 23360 25812 23394 26860
rect 23550 25812 23584 26860
rect 24756 25812 24790 26860
rect 24946 25812 24980 26860
rect 26152 25812 26186 26860
rect 26342 25812 26376 26860
rect 27548 25812 27582 26860
rect 27738 25812 27772 26860
rect 28944 25812 28978 26860
rect 29134 25812 29168 26860
rect 30340 25812 30374 26860
rect 30530 25812 30564 26860
rect 31736 25812 31770 26860
rect 31926 25812 31960 26860
rect 33132 25812 33166 26860
rect 33322 25812 33356 26860
rect 34528 25812 34562 26860
rect 34718 25812 34752 26860
rect 35924 25812 35958 26860
rect 36114 25812 36148 26860
rect 37320 25812 37354 26860
rect 37510 25812 37544 26860
rect 38716 25812 38750 26860
rect 38906 25812 38940 26860
rect 40112 25812 40146 26860
rect 40302 25812 40336 26860
rect 41508 25812 41542 26860
rect 41698 25812 41732 26860
rect 42904 25812 42938 26860
rect 43094 25812 43128 26860
rect 44300 25812 44334 26860
rect 44490 25812 44524 26860
rect 45696 25812 45730 26860
rect 45886 25812 45920 26860
rect 47092 25812 47126 26860
rect 47282 25812 47316 26860
rect 48488 25812 48522 26860
rect 48678 25812 48712 26860
rect 49884 25812 49918 26860
rect 50074 25812 50108 26860
rect 51280 25812 51314 26860
rect 9686 25716 9786 25750
rect 10634 25716 10734 25750
rect 11082 25716 11182 25750
rect 12030 25716 12130 25750
rect 12478 25716 12578 25750
rect 13426 25716 13526 25750
rect 13874 25716 13974 25750
rect 14822 25716 14922 25750
rect 15270 25716 15370 25750
rect 16218 25716 16318 25750
rect 16666 25716 16766 25750
rect 17614 25716 17714 25750
rect 18062 25716 18162 25750
rect 19010 25716 19110 25750
rect 19458 25716 19558 25750
rect 20406 25716 20506 25750
rect 20854 25716 20954 25750
rect 21802 25716 21902 25750
rect 22250 25716 22350 25750
rect 23198 25716 23298 25750
rect 23646 25716 23746 25750
rect 24594 25716 24694 25750
rect 25042 25716 25142 25750
rect 25990 25716 26090 25750
rect 26438 25716 26538 25750
rect 27386 25716 27486 25750
rect 27834 25716 27934 25750
rect 28782 25716 28882 25750
rect 29230 25716 29330 25750
rect 30178 25716 30278 25750
rect 30626 25716 30726 25750
rect 31574 25716 31674 25750
rect 32022 25716 32122 25750
rect 32970 25716 33070 25750
rect 33418 25716 33518 25750
rect 34366 25716 34466 25750
rect 34814 25716 34914 25750
rect 35762 25716 35862 25750
rect 36210 25716 36310 25750
rect 37158 25716 37258 25750
rect 37606 25716 37706 25750
rect 38554 25716 38654 25750
rect 39002 25716 39102 25750
rect 39950 25716 40050 25750
rect 40398 25716 40498 25750
rect 41346 25716 41446 25750
rect 41794 25716 41894 25750
rect 42742 25716 42842 25750
rect 43190 25716 43290 25750
rect 44138 25716 44238 25750
rect 44586 25716 44686 25750
rect 45534 25716 45634 25750
rect 45982 25716 46082 25750
rect 46930 25716 47030 25750
rect 47378 25716 47478 25750
rect 48326 25716 48426 25750
rect 48774 25716 48874 25750
rect 49722 25716 49822 25750
rect 50170 25716 50270 25750
rect 51118 25716 51218 25750
rect 51490 25602 51524 28466
rect 9476 25506 51428 25540
rect 3718 24054 4078 24414
rect -2944 18664 -2592 19016
rect 538 13412 604 13426
rect 360 13378 3630 13412
rect 538 13370 604 13378
rect 264 12074 298 13316
rect 3692 12074 3726 13316
rect 264 10098 298 11340
rect 3692 10098 3726 11340
rect 544 10036 3446 10038
rect 360 10002 3630 10036
<< metal1 >>
rect -1780 30854 7346 30864
rect -1780 30274 -1522 30854
rect 7242 30274 7346 30854
rect -1780 30264 7346 30274
rect -1780 30214 -1408 30264
rect -18962 30044 -2390 30046
rect -18962 30034 -2386 30044
rect -18962 29446 -2982 30034
rect -18962 28068 -18362 29446
rect -17410 29096 -17216 29102
rect -17792 28872 -17584 28880
rect -17792 28472 -17786 28872
rect -17590 28472 -17584 28872
rect -17792 28466 -17584 28472
rect -17410 28254 -17404 29096
rect -17222 28254 -17216 29096
rect -17410 28248 -17216 28254
rect -17184 28068 -16786 29446
rect -16004 29096 -15810 29102
rect -16386 28872 -16178 28880
rect -16386 28472 -16380 28872
rect -16184 28472 -16178 28872
rect -16386 28466 -16178 28472
rect -16004 28254 -15998 29096
rect -15816 28254 -15810 29096
rect -16004 28248 -15810 28254
rect -15778 28068 -15380 29446
rect -14598 29096 -14404 29102
rect -14980 28872 -14772 28880
rect -14980 28472 -14974 28872
rect -14778 28472 -14772 28872
rect -14980 28466 -14772 28472
rect -14598 28254 -14592 29096
rect -14410 28254 -14404 29096
rect -14598 28248 -14404 28254
rect -14372 28068 -13974 29446
rect -13192 29096 -12998 29102
rect -13574 28872 -13366 28880
rect -13574 28472 -13568 28872
rect -13372 28472 -13366 28872
rect -13574 28466 -13366 28472
rect -13192 28254 -13186 29096
rect -13004 28254 -12998 29096
rect -13192 28248 -12998 28254
rect -12966 28068 -12568 29446
rect -11786 29096 -11592 29102
rect -12168 28872 -11960 28880
rect -12168 28472 -12162 28872
rect -11966 28472 -11960 28872
rect -12168 28466 -11960 28472
rect -11786 28254 -11780 29096
rect -11598 28254 -11592 29096
rect -11786 28248 -11592 28254
rect -11560 28068 -11162 29446
rect -10380 29096 -10186 29102
rect -10762 28872 -10554 28880
rect -10762 28472 -10756 28872
rect -10560 28472 -10554 28872
rect -10762 28466 -10554 28472
rect -10380 28254 -10374 29096
rect -10192 28254 -10186 29096
rect -10380 28248 -10186 28254
rect -10154 28068 -9756 29446
rect -8974 29096 -8780 29102
rect -9356 28872 -9148 28880
rect -9356 28472 -9350 28872
rect -9154 28472 -9148 28872
rect -9356 28466 -9148 28472
rect -8974 28254 -8968 29096
rect -8786 28254 -8780 29096
rect -8974 28248 -8780 28254
rect -8748 28068 -8350 29446
rect -7568 29096 -7374 29102
rect -7950 28872 -7742 28880
rect -7950 28472 -7944 28872
rect -7748 28472 -7742 28872
rect -7950 28466 -7742 28472
rect -7568 28254 -7562 29096
rect -7380 28254 -7374 29096
rect -7568 28248 -7374 28254
rect -7342 28068 -6944 29446
rect -6162 29096 -5968 29102
rect -6544 28872 -6336 28880
rect -6544 28472 -6538 28872
rect -6342 28472 -6336 28872
rect -6544 28466 -6336 28472
rect -6162 28254 -6156 29096
rect -5974 28254 -5968 29096
rect -6162 28248 -5968 28254
rect -5936 28068 -5538 29446
rect -4362 29246 -3762 29446
rect -2992 29246 -2982 29446
rect -4756 29096 -4562 29102
rect -5138 28872 -4930 28880
rect -5138 28472 -5132 28872
rect -4936 28472 -4930 28872
rect -5138 28466 -4930 28472
rect -4756 28254 -4750 29096
rect -4568 28254 -4562 29096
rect -4756 28248 -4562 28254
rect -4362 28646 -2982 29246
rect -4362 28446 -3762 28646
rect -2992 28446 -2982 28646
rect -4362 28068 -2982 28446
rect -18962 27846 -2982 28068
rect -18962 27670 -3762 27846
rect -18962 26462 -18362 27670
rect -17410 27490 -17216 27496
rect -17792 27266 -17584 27274
rect -17792 26866 -17786 27266
rect -17590 26866 -17584 27266
rect -17792 26860 -17584 26866
rect -17410 26648 -17404 27490
rect -17222 26648 -17216 27490
rect -17410 26642 -17216 26648
rect -17184 26462 -16786 27670
rect -16004 27490 -15810 27496
rect -16386 27266 -16178 27274
rect -16386 26866 -16380 27266
rect -16184 26866 -16178 27266
rect -16386 26860 -16178 26866
rect -16004 26648 -15998 27490
rect -15816 26648 -15810 27490
rect -16004 26642 -15810 26648
rect -15778 26462 -15380 27670
rect -14598 27490 -14404 27496
rect -14980 27266 -14772 27274
rect -14980 26866 -14974 27266
rect -14778 26866 -14772 27266
rect -14980 26860 -14772 26866
rect -14598 26648 -14592 27490
rect -14410 26648 -14404 27490
rect -14598 26642 -14404 26648
rect -14372 26462 -13974 27670
rect -13192 27490 -12998 27496
rect -13574 27266 -13366 27274
rect -13574 26866 -13568 27266
rect -13372 26866 -13366 27266
rect -13574 26860 -13366 26866
rect -13192 26648 -13186 27490
rect -13004 26648 -12998 27490
rect -13192 26642 -12998 26648
rect -12966 26462 -12568 27670
rect -11786 27490 -11592 27496
rect -12168 27266 -11960 27274
rect -12168 26866 -12162 27266
rect -11966 26866 -11960 27266
rect -12168 26860 -11960 26866
rect -11786 26648 -11780 27490
rect -11598 26648 -11592 27490
rect -11786 26642 -11592 26648
rect -11560 26462 -11162 27670
rect -10380 27490 -10186 27496
rect -10762 27266 -10554 27274
rect -10762 26866 -10756 27266
rect -10560 26866 -10554 27266
rect -10762 26860 -10554 26866
rect -10380 26648 -10374 27490
rect -10192 26648 -10186 27490
rect -10380 26642 -10186 26648
rect -10154 26462 -9756 27670
rect -8974 27490 -8780 27496
rect -9356 27266 -9148 27274
rect -9356 26866 -9350 27266
rect -9154 26866 -9148 27266
rect -9356 26860 -9148 26866
rect -8974 26648 -8968 27490
rect -8786 26648 -8780 27490
rect -8974 26642 -8780 26648
rect -8748 26462 -8350 27670
rect -7568 27490 -7374 27496
rect -7950 27266 -7742 27274
rect -7950 26866 -7944 27266
rect -7748 26866 -7742 27266
rect -7950 26860 -7742 26866
rect -7568 26648 -7562 27490
rect -7380 26648 -7374 27490
rect -7568 26642 -7374 26648
rect -7342 26462 -6944 27670
rect -6162 27490 -5968 27496
rect -6544 27266 -6336 27274
rect -6544 26866 -6538 27266
rect -6342 26866 -6336 27266
rect -6544 26860 -6336 26866
rect -6162 26648 -6156 27490
rect -5974 26648 -5968 27490
rect -6162 26642 -5968 26648
rect -5936 26462 -5538 27670
rect -4362 27646 -3762 27670
rect -2992 27646 -2982 27846
rect -4756 27490 -4562 27496
rect -5138 27266 -4930 27274
rect -5138 26866 -5132 27266
rect -4936 26866 -4930 27266
rect -5138 26860 -4930 26866
rect -4756 26648 -4750 27490
rect -4568 26648 -4562 27490
rect -4756 26642 -4562 26648
rect -4362 27046 -2982 27646
rect -4362 26846 -3762 27046
rect -2992 26846 -2982 27046
rect -4362 26462 -2982 26846
rect -18962 26246 -2982 26462
rect -18962 26064 -3762 26246
rect -18962 24856 -18362 26064
rect -17410 25884 -17216 25890
rect -17792 25660 -17584 25668
rect -17792 25260 -17786 25660
rect -17590 25260 -17584 25660
rect -17792 25254 -17584 25260
rect -17410 25042 -17404 25884
rect -17222 25042 -17216 25884
rect -17410 25036 -17216 25042
rect -17184 24856 -16786 26064
rect -16004 25884 -15810 25890
rect -16386 25660 -16178 25668
rect -16386 25260 -16380 25660
rect -16184 25260 -16178 25660
rect -16386 25254 -16178 25260
rect -16004 25042 -15998 25884
rect -15816 25042 -15810 25884
rect -16004 25036 -15810 25042
rect -15778 24856 -15380 26064
rect -14598 25884 -14404 25890
rect -14980 25660 -14772 25668
rect -14980 25260 -14974 25660
rect -14778 25260 -14772 25660
rect -14980 25254 -14772 25260
rect -14598 25042 -14592 25884
rect -14410 25042 -14404 25884
rect -14598 25036 -14404 25042
rect -14372 24856 -13974 26064
rect -13192 25884 -12998 25890
rect -13574 25660 -13366 25668
rect -13574 25260 -13568 25660
rect -13372 25260 -13366 25660
rect -13574 25254 -13366 25260
rect -13192 25042 -13186 25884
rect -13004 25042 -12998 25884
rect -13192 25036 -12998 25042
rect -12966 24856 -12568 26064
rect -11786 25884 -11592 25890
rect -12168 25660 -11960 25668
rect -12168 25260 -12162 25660
rect -11966 25260 -11960 25660
rect -12168 25254 -11960 25260
rect -11786 25042 -11780 25884
rect -11598 25042 -11592 25884
rect -11786 25036 -11592 25042
rect -11560 24856 -11162 26064
rect -10380 25884 -10186 25890
rect -10762 25660 -10554 25668
rect -10762 25260 -10756 25660
rect -10560 25260 -10554 25660
rect -10762 25254 -10554 25260
rect -10380 25042 -10374 25884
rect -10192 25042 -10186 25884
rect -10380 25036 -10186 25042
rect -10154 24856 -9756 26064
rect -8974 25884 -8780 25890
rect -9356 25660 -9148 25668
rect -9356 25260 -9350 25660
rect -9154 25260 -9148 25660
rect -9356 25254 -9148 25260
rect -8974 25042 -8968 25884
rect -8786 25042 -8780 25884
rect -8974 25036 -8780 25042
rect -8748 24856 -8350 26064
rect -7568 25884 -7374 25890
rect -7950 25660 -7742 25668
rect -7950 25260 -7944 25660
rect -7748 25260 -7742 25660
rect -7950 25254 -7742 25260
rect -7568 25042 -7562 25884
rect -7380 25042 -7374 25884
rect -7568 25036 -7374 25042
rect -7342 24856 -6944 26064
rect -6162 25884 -5968 25890
rect -6544 25660 -6336 25668
rect -6544 25260 -6538 25660
rect -6342 25260 -6336 25660
rect -6544 25254 -6336 25260
rect -6162 25042 -6156 25884
rect -5974 25042 -5968 25884
rect -6162 25036 -5968 25042
rect -5936 24856 -5538 26064
rect -4362 26046 -3762 26064
rect -2992 26046 -2982 26246
rect -4756 25884 -4562 25890
rect -5138 25660 -4930 25668
rect -5138 25260 -5132 25660
rect -4936 25260 -4930 25660
rect -5138 25254 -4930 25260
rect -4756 25042 -4750 25884
rect -4568 25042 -4562 25884
rect -4756 25036 -4562 25042
rect -4362 25446 -2982 26046
rect -4362 25246 -3762 25446
rect -2992 25246 -2982 25446
rect -4362 24856 -2982 25246
rect -18962 24656 -2982 24856
rect -2396 24656 -2386 30034
rect -18962 24646 -2386 24656
rect -1780 29166 -1454 30214
rect -1420 29166 -1408 30214
rect -260 30214 -12 30264
rect -1234 30080 -434 30090
rect -1234 29300 -1224 30080
rect -444 29300 -434 30080
rect -1234 29290 -434 29300
rect -1780 29116 -1408 29166
rect -260 29166 -248 30214
rect -214 29166 -58 30214
rect -24 29166 -12 30214
rect 1136 30214 1384 30264
rect 162 30080 962 30090
rect 162 29300 172 30080
rect 952 29300 962 30080
rect 162 29290 962 29300
rect -260 29116 -12 29166
rect 1136 29166 1148 30214
rect 1182 29166 1338 30214
rect 1372 29166 1384 30214
rect 2532 30214 2780 30264
rect 1558 30080 2358 30090
rect 1558 29300 1568 30080
rect 2348 29300 2358 30080
rect 1558 29290 2358 29300
rect 1136 29116 1384 29166
rect 2532 29166 2544 30214
rect 2578 29166 2734 30214
rect 2768 29166 2780 30214
rect 3928 30214 4298 30264
rect 2954 30080 3754 30090
rect 2954 29300 2964 30080
rect 3744 29300 3754 30080
rect 2954 29290 3754 29300
rect 2532 29116 2780 29166
rect 3928 29166 3940 30214
rect 3974 29166 4298 30214
rect 3928 29116 4298 29166
rect -1780 29106 4298 29116
rect -1780 28878 -1696 29106
rect -1368 29104 -300 29106
rect -1368 29070 -1358 29104
rect -310 29070 -300 29104
rect -1368 28914 -300 29070
rect -1368 28880 -1358 28914
rect -310 28880 -300 28914
rect -1368 28878 -300 28880
rect 28 29104 1096 29106
rect 28 29070 38 29104
rect 1086 29070 1096 29104
rect 28 28914 1096 29070
rect 28 28880 38 28914
rect 1086 28880 1096 28914
rect 28 28878 1096 28880
rect 1424 29104 2492 29106
rect 1424 29070 1434 29104
rect 2482 29070 2492 29104
rect 1424 28914 2492 29070
rect 1424 28880 1434 28914
rect 2482 28880 2492 28914
rect 1424 28878 2492 28880
rect 2820 29104 3888 29106
rect 2820 29070 2830 29104
rect 3878 29070 3888 29104
rect 2820 28914 3888 29070
rect 2820 28880 2830 28914
rect 3878 28880 3888 28914
rect 2820 28878 3888 28880
rect 4216 28878 4298 29106
rect -1780 28868 4298 28878
rect -1780 28818 -1408 28868
rect -1780 27770 -1454 28818
rect -1420 27770 -1408 28818
rect -260 28818 -12 28868
rect -1234 28684 -434 28694
rect -1234 27904 -1224 28684
rect -444 27904 -434 28684
rect -1234 27894 -434 27904
rect -1780 27720 -1408 27770
rect -260 27770 -248 28818
rect -214 27770 -58 28818
rect -24 27770 -12 28818
rect 1136 28818 1384 28868
rect 162 28684 962 28694
rect 162 27904 172 28684
rect 952 27904 962 28684
rect 162 27894 962 27904
rect -260 27720 -12 27770
rect 1136 27770 1148 28818
rect 1182 27770 1338 28818
rect 1372 27770 1384 28818
rect 2532 28818 2780 28868
rect 1558 28684 2358 28694
rect 1558 27904 1568 28684
rect 2348 27904 2358 28684
rect 1558 27894 2358 27904
rect 1136 27720 1384 27770
rect 2532 27770 2544 28818
rect 2578 27770 2734 28818
rect 2768 27770 2780 28818
rect 3928 28818 4298 28868
rect 2954 28684 3754 28694
rect 2954 27904 2964 28684
rect 3744 27904 3754 28684
rect 2954 27894 3754 27904
rect 2532 27720 2780 27770
rect 3928 27770 3940 28818
rect 3974 27770 4298 28818
rect 3928 27720 4298 27770
rect -1780 27710 4298 27720
rect -1780 27482 -1696 27710
rect -1368 27708 -300 27710
rect -1368 27674 -1358 27708
rect -310 27674 -300 27708
rect -1368 27518 -300 27674
rect -1368 27484 -1358 27518
rect -310 27484 -300 27518
rect -1368 27482 -300 27484
rect 28 27708 1096 27710
rect 28 27674 38 27708
rect 1086 27674 1096 27708
rect 28 27518 1096 27674
rect 28 27484 38 27518
rect 1086 27484 1096 27518
rect 28 27482 1096 27484
rect 1424 27708 2492 27710
rect 1424 27674 1434 27708
rect 2482 27674 2492 27708
rect 1424 27518 2492 27674
rect 1424 27484 1434 27518
rect 2482 27484 2492 27518
rect 1424 27482 2492 27484
rect 2820 27708 3888 27710
rect 2820 27674 2830 27708
rect 3878 27674 3888 27708
rect 2820 27518 3888 27674
rect 2820 27484 2830 27518
rect 3878 27484 3888 27518
rect 2820 27482 3888 27484
rect 4216 27482 4298 27710
rect -1780 27472 4298 27482
rect -1780 27422 -1408 27472
rect -1780 26374 -1454 27422
rect -1420 26374 -1408 27422
rect -260 27422 -12 27472
rect -1234 27288 -434 27298
rect -1234 26508 -1224 27288
rect -444 26508 -434 27288
rect -1234 26498 -434 26508
rect -1780 26324 -1408 26374
rect -260 26374 -248 27422
rect -214 26374 -58 27422
rect -24 26374 -12 27422
rect 1136 27422 1384 27472
rect 162 27288 962 27298
rect 162 26508 172 27288
rect 952 26508 962 27288
rect 162 26498 962 26508
rect -260 26324 -12 26374
rect 1136 26374 1148 27422
rect 1182 26374 1338 27422
rect 1372 26374 1384 27422
rect 2532 27422 2780 27472
rect 1558 27288 2358 27298
rect 1558 26508 1568 27288
rect 2348 26508 2358 27288
rect 1558 26498 2358 26508
rect 1136 26324 1384 26374
rect 2532 26374 2544 27422
rect 2578 26374 2734 27422
rect 2768 26374 2780 27422
rect 3928 27422 4298 27472
rect 2954 27288 3754 27298
rect 2954 26508 2964 27288
rect 3744 26508 3754 27288
rect 2954 26498 3754 26508
rect 2532 26324 2780 26374
rect 3928 26374 3940 27422
rect 3974 26374 4298 27422
rect 3928 26324 4298 26374
rect -1780 26314 4298 26324
rect -1780 26086 -1696 26314
rect -1368 26312 -300 26314
rect -1368 26278 -1358 26312
rect -310 26278 -300 26312
rect -1368 26122 -300 26278
rect -1368 26088 -1358 26122
rect -310 26088 -300 26122
rect -1368 26086 -300 26088
rect 28 26312 1096 26314
rect 28 26278 38 26312
rect 1086 26278 1096 26312
rect 28 26122 1096 26278
rect 28 26088 38 26122
rect 1086 26088 1096 26122
rect 28 26086 1096 26088
rect 1424 26312 2492 26314
rect 1424 26278 1434 26312
rect 2482 26278 2492 26312
rect 1424 26122 2492 26278
rect 1424 26088 1434 26122
rect 2482 26088 2492 26122
rect 1424 26086 2492 26088
rect 2820 26312 3888 26314
rect 2820 26278 2830 26312
rect 3878 26278 3888 26312
rect 2820 26122 3888 26278
rect 2820 26088 2830 26122
rect 3878 26088 3888 26122
rect 2820 26086 3888 26088
rect 4216 26086 4298 26314
rect -1780 26076 4298 26086
rect -1780 26026 -1408 26076
rect -1780 24978 -1454 26026
rect -1420 24978 -1408 26026
rect -260 26026 -12 26076
rect -1234 25892 -434 25902
rect -1234 25112 -1224 25892
rect -444 25112 -434 25892
rect -1234 25102 -434 25112
rect -1780 24928 -1408 24978
rect -260 24978 -248 26026
rect -214 24978 -58 26026
rect -24 24978 -12 26026
rect 1136 26026 1384 26076
rect 162 25892 962 25902
rect 162 25112 172 25892
rect 952 25112 962 25892
rect 162 25102 962 25112
rect -260 24928 -12 24978
rect 1136 24978 1148 26026
rect 1182 24978 1338 26026
rect 1372 24978 1384 26026
rect 2532 26026 2780 26076
rect 1558 25892 2358 25902
rect 1558 25112 1568 25892
rect 2348 25112 2358 25892
rect 1558 25102 2358 25112
rect 1136 24928 1384 24978
rect 2532 24978 2544 26026
rect 2578 24978 2734 26026
rect 2768 24978 2780 26026
rect 3928 26026 4298 26076
rect 2954 25892 3754 25902
rect 2954 25112 2964 25892
rect 3744 25112 3754 25892
rect 2954 25102 3754 25112
rect 2532 24928 2780 24978
rect 3928 24978 3940 26026
rect 3974 24978 4298 26026
rect 9368 28562 51536 28574
rect 9368 28528 9476 28562
rect 51428 28528 51536 28562
rect 9368 28516 51536 28528
rect 9368 28466 9426 28516
rect 9368 25602 9380 28466
rect 9414 25602 9426 28466
rect 51478 28466 51536 28516
rect 9512 28352 51392 28430
rect 9512 28318 9686 28352
rect 10734 28318 11082 28352
rect 12130 28318 12478 28352
rect 13526 28318 13874 28352
rect 14922 28318 15270 28352
rect 16318 28318 16666 28352
rect 17714 28318 18062 28352
rect 19110 28318 19458 28352
rect 20506 28318 20854 28352
rect 21902 28318 22250 28352
rect 23298 28318 23646 28352
rect 24694 28318 25042 28352
rect 26090 28318 26438 28352
rect 27486 28318 27834 28352
rect 28882 28318 29230 28352
rect 30278 28318 30626 28352
rect 31674 28318 32022 28352
rect 33070 28318 33418 28352
rect 34466 28318 34814 28352
rect 35862 28318 36210 28352
rect 37258 28318 37606 28352
rect 38654 28318 39002 28352
rect 40050 28318 40398 28352
rect 41446 28318 41794 28352
rect 42842 28318 43190 28352
rect 44238 28318 44586 28352
rect 45634 28318 45982 28352
rect 47030 28318 47378 28352
rect 48426 28318 48774 28352
rect 49822 28318 50170 28352
rect 51218 28318 51392 28352
rect 9512 28306 51392 28318
rect 9512 28256 9636 28306
rect 9512 27208 9590 28256
rect 9624 27208 9636 28256
rect 10784 28256 11032 28306
rect 9710 28122 10710 28226
rect 9710 27342 9820 28122
rect 10600 27342 10710 28122
rect 9710 27238 10710 27342
rect 9512 27158 9636 27208
rect 10784 27158 10796 28256
rect 9512 27146 9792 27158
rect 9512 27112 9686 27146
rect 9786 27112 9792 27146
rect 9512 27100 9792 27112
rect 10628 27146 10796 27158
rect 10628 27112 10634 27146
rect 10734 27112 10796 27146
rect 10628 27100 10796 27112
rect 9512 26968 9636 27100
rect 10784 26968 10796 27100
rect 9512 26956 9792 26968
rect 9512 26922 9686 26956
rect 9786 26922 9792 26956
rect 9512 26910 9792 26922
rect 10628 26956 10796 26968
rect 10628 26922 10634 26956
rect 10734 26922 10796 26956
rect 10628 26910 10796 26922
rect 9512 26860 9636 26910
rect 9512 25812 9590 26860
rect 9624 25812 9636 26860
rect 9710 26726 10710 26830
rect 9710 25946 9820 26726
rect 10600 25946 10710 26726
rect 9710 25842 10710 25946
rect 9512 25762 9636 25812
rect 10784 25762 10796 26910
rect 11020 27158 11032 28256
rect 12180 28256 12428 28306
rect 11106 28122 12106 28226
rect 11106 27342 11216 28122
rect 11996 27342 12106 28122
rect 11106 27238 12106 27342
rect 12180 27158 12192 28256
rect 11020 27146 11188 27158
rect 11020 27112 11082 27146
rect 11182 27112 11188 27146
rect 11020 27100 11188 27112
rect 12024 27146 12192 27158
rect 12024 27112 12030 27146
rect 12130 27112 12192 27146
rect 12024 27100 12192 27112
rect 11020 26968 11032 27100
rect 12180 26968 12192 27100
rect 11020 26956 11188 26968
rect 11020 26922 11082 26956
rect 11182 26922 11188 26956
rect 11020 26910 11188 26922
rect 12024 26956 12192 26968
rect 12024 26922 12030 26956
rect 12130 26922 12192 26956
rect 12024 26910 12192 26922
rect 9512 25750 9792 25762
rect 9512 25716 9686 25750
rect 9786 25716 9792 25750
rect 9512 25704 9792 25716
rect 10628 25750 10796 25762
rect 10628 25716 10634 25750
rect 10734 25716 10796 25750
rect 11020 25762 11032 26910
rect 11106 26726 12106 26830
rect 11106 25946 11216 26726
rect 11996 25946 12106 26726
rect 11106 25842 12106 25946
rect 12180 25762 12192 26910
rect 12416 27158 12428 28256
rect 13576 28256 13824 28306
rect 12510 28122 13502 28226
rect 12510 27342 12612 28122
rect 13392 27342 13502 28122
rect 12510 27238 13502 27342
rect 13576 27158 13588 28256
rect 12416 27146 12584 27158
rect 12416 27112 12478 27146
rect 12578 27112 12584 27146
rect 12416 27100 12584 27112
rect 13420 27146 13588 27158
rect 13420 27112 13426 27146
rect 13526 27112 13588 27146
rect 13420 27100 13588 27112
rect 12416 26968 12428 27100
rect 13576 26968 13588 27100
rect 12416 26956 12584 26968
rect 12416 26922 12478 26956
rect 12578 26922 12584 26956
rect 12416 26910 12584 26922
rect 13420 26956 13588 26968
rect 13420 26922 13426 26956
rect 13526 26922 13588 26956
rect 13420 26910 13588 26922
rect 11020 25750 11188 25762
rect 11020 25716 11082 25750
rect 11182 25716 11188 25750
rect 10628 25704 11188 25716
rect 12024 25750 12192 25762
rect 12024 25716 12030 25750
rect 12130 25716 12192 25750
rect 12416 25762 12428 26910
rect 12510 26726 13502 26830
rect 12510 25946 12612 26726
rect 13392 25946 13502 26726
rect 12510 25842 13502 25946
rect 13576 25762 13588 26910
rect 13812 27158 13824 28256
rect 14972 28256 15220 28306
rect 13898 28122 14898 28226
rect 13898 27342 14008 28122
rect 14788 27342 14898 28122
rect 13898 27238 14898 27342
rect 14972 27158 14984 28256
rect 13812 27146 13980 27158
rect 13812 27112 13874 27146
rect 13974 27112 13980 27146
rect 13812 27100 13980 27112
rect 14816 27146 14984 27158
rect 14816 27112 14822 27146
rect 14922 27112 14984 27146
rect 14816 27100 14984 27112
rect 13812 26968 13824 27100
rect 14972 26968 14984 27100
rect 13812 26956 13980 26968
rect 13812 26922 13874 26956
rect 13974 26922 13980 26956
rect 13812 26910 13980 26922
rect 14816 26956 14984 26968
rect 14816 26922 14822 26956
rect 14922 26922 14984 26956
rect 14816 26910 14984 26922
rect 12416 25750 12584 25762
rect 12416 25716 12478 25750
rect 12578 25716 12584 25750
rect 12024 25704 12584 25716
rect 13420 25750 13588 25762
rect 13420 25716 13426 25750
rect 13526 25716 13588 25750
rect 13812 25762 13824 26910
rect 13898 26726 14898 26830
rect 13898 25946 14008 26726
rect 14788 25946 14898 26726
rect 13898 25842 14898 25946
rect 14972 25762 14984 26910
rect 15208 27158 15220 28256
rect 16368 28256 16616 28306
rect 15294 28122 16294 28226
rect 15294 27342 15404 28122
rect 16184 27342 16294 28122
rect 15294 27238 16294 27342
rect 16368 27158 16380 28256
rect 15208 27146 15376 27158
rect 15208 27112 15270 27146
rect 15370 27112 15376 27146
rect 15208 27100 15376 27112
rect 16212 27146 16380 27158
rect 16212 27112 16218 27146
rect 16318 27112 16380 27146
rect 16212 27100 16380 27112
rect 15208 26968 15220 27100
rect 16368 26968 16380 27100
rect 15208 26956 15376 26968
rect 15208 26922 15270 26956
rect 15370 26922 15376 26956
rect 15208 26910 15376 26922
rect 16212 26956 16380 26968
rect 16212 26922 16218 26956
rect 16318 26922 16380 26956
rect 16212 26910 16380 26922
rect 13812 25750 13980 25762
rect 13812 25716 13874 25750
rect 13974 25716 13980 25750
rect 13420 25704 13980 25716
rect 14816 25750 14984 25762
rect 14816 25716 14822 25750
rect 14922 25716 14984 25750
rect 15208 25762 15220 26910
rect 15294 26726 16294 26830
rect 15294 25946 15404 26726
rect 16184 25946 16294 26726
rect 15294 25842 16294 25946
rect 16368 25762 16380 26910
rect 16604 27158 16616 28256
rect 17764 28256 18012 28306
rect 16690 28122 17690 28226
rect 16690 27342 16800 28122
rect 17580 27342 17690 28122
rect 16690 27238 17690 27342
rect 17764 27158 17776 28256
rect 16604 27146 16772 27158
rect 16604 27112 16666 27146
rect 16766 27112 16772 27146
rect 16604 27100 16772 27112
rect 17608 27146 17776 27158
rect 17608 27112 17614 27146
rect 17714 27112 17776 27146
rect 17608 27100 17776 27112
rect 16604 26968 16616 27100
rect 17764 26968 17776 27100
rect 16604 26956 16772 26968
rect 16604 26922 16666 26956
rect 16766 26922 16772 26956
rect 16604 26910 16772 26922
rect 17608 26956 17776 26968
rect 17608 26922 17614 26956
rect 17714 26922 17776 26956
rect 17608 26910 17776 26922
rect 15208 25750 15376 25762
rect 15208 25716 15270 25750
rect 15370 25716 15376 25750
rect 14816 25704 15376 25716
rect 16212 25750 16380 25762
rect 16212 25716 16218 25750
rect 16318 25716 16380 25750
rect 16604 25762 16616 26910
rect 16690 26726 17690 26830
rect 16690 25946 16800 26726
rect 17580 25946 17690 26726
rect 16690 25842 17690 25946
rect 17764 25762 17776 26910
rect 18000 27158 18012 28256
rect 19160 28256 19408 28306
rect 18086 28122 19086 28226
rect 18086 27342 18196 28122
rect 18976 27342 19086 28122
rect 18086 27238 19086 27342
rect 19160 27158 19172 28256
rect 18000 27146 18168 27158
rect 18000 27112 18062 27146
rect 18162 27112 18168 27146
rect 18000 27100 18168 27112
rect 19004 27146 19172 27158
rect 19004 27112 19010 27146
rect 19110 27112 19172 27146
rect 19004 27100 19172 27112
rect 18000 26968 18012 27100
rect 19160 26968 19172 27100
rect 18000 26956 18168 26968
rect 18000 26922 18062 26956
rect 18162 26922 18168 26956
rect 18000 26910 18168 26922
rect 19004 26956 19172 26968
rect 19004 26922 19010 26956
rect 19110 26922 19172 26956
rect 19004 26910 19172 26922
rect 16604 25750 16772 25762
rect 16604 25716 16666 25750
rect 16766 25716 16772 25750
rect 16212 25704 16772 25716
rect 17608 25750 17776 25762
rect 17608 25716 17614 25750
rect 17714 25716 17776 25750
rect 18000 25762 18012 26910
rect 18086 26726 19086 26830
rect 18086 25946 18196 26726
rect 18976 25946 19086 26726
rect 18086 25842 19086 25946
rect 19160 25762 19172 26910
rect 19396 27158 19408 28256
rect 20556 28256 20804 28306
rect 19482 28122 20482 28226
rect 19482 27342 19592 28122
rect 20372 27342 20482 28122
rect 19482 27238 20482 27342
rect 20556 27158 20568 28256
rect 19396 27146 19564 27158
rect 19396 27112 19458 27146
rect 19558 27112 19564 27146
rect 19396 27100 19564 27112
rect 20400 27146 20568 27158
rect 20400 27112 20406 27146
rect 20506 27112 20568 27146
rect 20400 27100 20568 27112
rect 19396 26968 19408 27100
rect 20556 26968 20568 27100
rect 19396 26956 19564 26968
rect 19396 26922 19458 26956
rect 19558 26922 19564 26956
rect 19396 26910 19564 26922
rect 20400 26956 20568 26968
rect 20400 26922 20406 26956
rect 20506 26922 20568 26956
rect 20400 26910 20568 26922
rect 18000 25750 18168 25762
rect 18000 25716 18062 25750
rect 18162 25716 18168 25750
rect 17608 25704 18168 25716
rect 19004 25750 19172 25762
rect 19004 25716 19010 25750
rect 19110 25716 19172 25750
rect 19396 25762 19408 26910
rect 19482 26726 20482 26830
rect 19482 25946 19592 26726
rect 20372 25946 20482 26726
rect 19482 25842 20482 25946
rect 20556 25762 20568 26910
rect 20792 27158 20804 28256
rect 21952 28256 22200 28306
rect 20878 28122 21878 28226
rect 20878 27342 20988 28122
rect 21768 27342 21878 28122
rect 20878 27238 21878 27342
rect 21952 27158 21964 28256
rect 20792 27146 20960 27158
rect 20792 27112 20854 27146
rect 20954 27112 20960 27146
rect 20792 27100 20960 27112
rect 21796 27146 21964 27158
rect 21796 27112 21802 27146
rect 21902 27112 21964 27146
rect 21796 27100 21964 27112
rect 20792 26968 20804 27100
rect 21952 26968 21964 27100
rect 20792 26956 20960 26968
rect 20792 26922 20854 26956
rect 20954 26922 20960 26956
rect 20792 26910 20960 26922
rect 21796 26956 21964 26968
rect 21796 26922 21802 26956
rect 21902 26922 21964 26956
rect 21796 26910 21964 26922
rect 19396 25750 19564 25762
rect 19396 25716 19458 25750
rect 19558 25716 19564 25750
rect 19004 25704 19564 25716
rect 20400 25750 20568 25762
rect 20400 25716 20406 25750
rect 20506 25716 20568 25750
rect 20792 25762 20804 26910
rect 20878 26726 21878 26830
rect 20878 25946 20988 26726
rect 21768 25946 21878 26726
rect 20878 25842 21878 25946
rect 21952 25762 21964 26910
rect 22188 27158 22200 28256
rect 23348 28256 23596 28306
rect 22274 28122 23274 28226
rect 22274 27342 22384 28122
rect 23164 27342 23274 28122
rect 22274 27238 23274 27342
rect 23348 27158 23360 28256
rect 22188 27146 22356 27158
rect 22188 27112 22250 27146
rect 22350 27112 22356 27146
rect 22188 27100 22356 27112
rect 23192 27146 23360 27158
rect 23192 27112 23198 27146
rect 23298 27112 23360 27146
rect 23192 27100 23360 27112
rect 22188 26968 22200 27100
rect 23348 26968 23360 27100
rect 22188 26956 22356 26968
rect 22188 26922 22250 26956
rect 22350 26922 22356 26956
rect 22188 26910 22356 26922
rect 23192 26956 23360 26968
rect 23192 26922 23198 26956
rect 23298 26922 23360 26956
rect 23192 26910 23360 26922
rect 20792 25750 20960 25762
rect 20792 25716 20854 25750
rect 20954 25716 20960 25750
rect 20400 25704 20960 25716
rect 21796 25750 21964 25762
rect 21796 25716 21802 25750
rect 21902 25716 21964 25750
rect 22188 25762 22200 26910
rect 22274 26726 23274 26830
rect 22274 25946 22384 26726
rect 23164 25946 23274 26726
rect 22274 25842 23274 25946
rect 23348 25762 23360 26910
rect 23584 27158 23596 28256
rect 24744 28256 24992 28306
rect 23670 28122 24670 28226
rect 23670 27342 23780 28122
rect 24560 27342 24670 28122
rect 23670 27238 24670 27342
rect 24744 27158 24756 28256
rect 23584 27146 23752 27158
rect 23584 27112 23646 27146
rect 23746 27112 23752 27146
rect 23584 27100 23752 27112
rect 24588 27146 24756 27158
rect 24588 27112 24594 27146
rect 24694 27112 24756 27146
rect 24588 27100 24756 27112
rect 23584 26968 23596 27100
rect 24744 26968 24756 27100
rect 23584 26956 23752 26968
rect 23584 26922 23646 26956
rect 23746 26922 23752 26956
rect 23584 26910 23752 26922
rect 24588 26956 24756 26968
rect 24588 26922 24594 26956
rect 24694 26922 24756 26956
rect 24588 26910 24756 26922
rect 22188 25750 22356 25762
rect 22188 25716 22250 25750
rect 22350 25716 22356 25750
rect 21796 25704 22356 25716
rect 23192 25750 23360 25762
rect 23192 25716 23198 25750
rect 23298 25716 23360 25750
rect 23584 25762 23596 26910
rect 23670 26726 24670 26830
rect 23670 25946 23780 26726
rect 24560 25946 24670 26726
rect 23670 25842 24670 25946
rect 24744 25762 24756 26910
rect 24980 27158 24992 28256
rect 26140 28256 26388 28306
rect 25066 28122 26066 28226
rect 25066 27342 25176 28122
rect 25956 27342 26066 28122
rect 25066 27238 26066 27342
rect 26140 27158 26152 28256
rect 24980 27146 25148 27158
rect 24980 27112 25042 27146
rect 25142 27112 25148 27146
rect 24980 27100 25148 27112
rect 25984 27146 26152 27158
rect 25984 27112 25990 27146
rect 26090 27112 26152 27146
rect 25984 27100 26152 27112
rect 24980 26968 24992 27100
rect 26140 26968 26152 27100
rect 24980 26956 25148 26968
rect 24980 26922 25042 26956
rect 25142 26922 25148 26956
rect 24980 26910 25148 26922
rect 25984 26956 26152 26968
rect 25984 26922 25990 26956
rect 26090 26922 26152 26956
rect 25984 26910 26152 26922
rect 23584 25750 23752 25762
rect 23584 25716 23646 25750
rect 23746 25716 23752 25750
rect 23192 25704 23752 25716
rect 24588 25750 24756 25762
rect 24588 25716 24594 25750
rect 24694 25716 24756 25750
rect 24980 25762 24992 26910
rect 25066 26726 26066 26830
rect 25066 25946 25176 26726
rect 25956 25946 26066 26726
rect 25066 25842 26066 25946
rect 26140 25762 26152 26910
rect 26376 27158 26388 28256
rect 27536 28256 27784 28306
rect 26462 28122 27462 28226
rect 26462 27342 26572 28122
rect 27352 27342 27462 28122
rect 26462 27238 27462 27342
rect 27536 27158 27548 28256
rect 26376 27146 26544 27158
rect 26376 27112 26438 27146
rect 26538 27112 26544 27146
rect 26376 27100 26544 27112
rect 27380 27146 27548 27158
rect 27380 27112 27386 27146
rect 27486 27112 27548 27146
rect 27380 27100 27548 27112
rect 26376 26968 26388 27100
rect 27536 26968 27548 27100
rect 26376 26956 26544 26968
rect 26376 26922 26438 26956
rect 26538 26922 26544 26956
rect 26376 26910 26544 26922
rect 27380 26956 27548 26968
rect 27380 26922 27386 26956
rect 27486 26922 27548 26956
rect 27380 26910 27548 26922
rect 24980 25750 25148 25762
rect 24980 25716 25042 25750
rect 25142 25716 25148 25750
rect 24588 25704 25148 25716
rect 25984 25750 26152 25762
rect 25984 25716 25990 25750
rect 26090 25716 26152 25750
rect 26376 25762 26388 26910
rect 26462 26726 27462 26830
rect 26462 25946 26572 26726
rect 27352 25946 27462 26726
rect 26462 25842 27462 25946
rect 27536 25762 27548 26910
rect 27772 27158 27784 28256
rect 28932 28256 29180 28306
rect 27858 28122 28858 28226
rect 27858 27342 27968 28122
rect 28748 27342 28858 28122
rect 27858 27238 28858 27342
rect 28932 27158 28944 28256
rect 27772 27146 27940 27158
rect 27772 27112 27834 27146
rect 27934 27112 27940 27146
rect 27772 27100 27940 27112
rect 28776 27146 28944 27158
rect 28776 27112 28782 27146
rect 28882 27112 28944 27146
rect 28776 27100 28944 27112
rect 27772 26968 27784 27100
rect 28932 26968 28944 27100
rect 27772 26956 27940 26968
rect 27772 26922 27834 26956
rect 27934 26922 27940 26956
rect 27772 26910 27940 26922
rect 28776 26956 28944 26968
rect 28776 26922 28782 26956
rect 28882 26922 28944 26956
rect 28776 26910 28944 26922
rect 26376 25750 26544 25762
rect 26376 25716 26438 25750
rect 26538 25716 26544 25750
rect 25984 25704 26544 25716
rect 27380 25750 27548 25762
rect 27380 25716 27386 25750
rect 27486 25716 27548 25750
rect 27772 25762 27784 26910
rect 27858 26726 28858 26830
rect 27858 25946 27968 26726
rect 28748 25946 28858 26726
rect 27858 25842 28858 25946
rect 28932 25762 28944 26910
rect 29168 27158 29180 28256
rect 30328 28256 30576 28306
rect 29252 28122 30254 28226
rect 29252 27342 29362 28122
rect 30144 27342 30254 28122
rect 29252 27238 30254 27342
rect 30328 27158 30340 28256
rect 29168 27146 29336 27158
rect 29168 27112 29230 27146
rect 29330 27112 29336 27146
rect 29168 27100 29336 27112
rect 30172 27146 30340 27158
rect 30172 27112 30178 27146
rect 30278 27112 30340 27146
rect 30172 27100 30340 27112
rect 29168 26968 29180 27100
rect 30328 26968 30340 27100
rect 29168 26956 29336 26968
rect 29168 26922 29230 26956
rect 29330 26922 29336 26956
rect 29168 26910 29336 26922
rect 30172 26956 30340 26968
rect 30172 26922 30178 26956
rect 30278 26922 30340 26956
rect 30172 26910 30340 26922
rect 27772 25750 27940 25762
rect 27772 25716 27834 25750
rect 27934 25716 27940 25750
rect 27380 25704 27940 25716
rect 28776 25750 28944 25762
rect 28776 25716 28782 25750
rect 28882 25716 28944 25750
rect 29168 25762 29180 26910
rect 29252 26726 30254 26830
rect 29252 25946 29362 26726
rect 30144 25946 30254 26726
rect 29252 25842 30254 25946
rect 30328 25762 30340 26910
rect 30564 27158 30576 28256
rect 31724 28256 31972 28306
rect 30650 28122 31650 28226
rect 30650 27342 30760 28122
rect 31540 27342 31650 28122
rect 30650 27238 31650 27342
rect 31724 27158 31736 28256
rect 30564 27146 30732 27158
rect 30564 27112 30626 27146
rect 30726 27112 30732 27146
rect 30564 27100 30732 27112
rect 31568 27146 31736 27158
rect 31568 27112 31574 27146
rect 31674 27112 31736 27146
rect 31568 27100 31736 27112
rect 30564 26968 30576 27100
rect 31724 26968 31736 27100
rect 30564 26956 30732 26968
rect 30564 26922 30626 26956
rect 30726 26922 30732 26956
rect 30564 26910 30732 26922
rect 31568 26956 31736 26968
rect 31568 26922 31574 26956
rect 31674 26922 31736 26956
rect 31568 26910 31736 26922
rect 29168 25750 29336 25762
rect 29168 25716 29230 25750
rect 29330 25716 29336 25750
rect 28776 25704 29336 25716
rect 30172 25750 30340 25762
rect 30172 25716 30178 25750
rect 30278 25716 30340 25750
rect 30564 25762 30576 26910
rect 30650 26726 31650 26830
rect 30650 25946 30760 26726
rect 31540 25946 31650 26726
rect 30650 25842 31650 25946
rect 31724 25762 31736 26910
rect 31960 27158 31972 28256
rect 33120 28256 33368 28306
rect 32046 28122 33046 28226
rect 32046 27342 32156 28122
rect 32936 27342 33046 28122
rect 32046 27238 33046 27342
rect 33120 27158 33132 28256
rect 31960 27146 32128 27158
rect 31960 27112 32022 27146
rect 32122 27112 32128 27146
rect 31960 27100 32128 27112
rect 32964 27146 33132 27158
rect 32964 27112 32970 27146
rect 33070 27112 33132 27146
rect 32964 27100 33132 27112
rect 31960 26968 31972 27100
rect 33120 26968 33132 27100
rect 31960 26956 32128 26968
rect 31960 26922 32022 26956
rect 32122 26922 32128 26956
rect 31960 26910 32128 26922
rect 32964 26956 33132 26968
rect 32964 26922 32970 26956
rect 33070 26922 33132 26956
rect 32964 26910 33132 26922
rect 30564 25750 30732 25762
rect 30564 25716 30626 25750
rect 30726 25716 30732 25750
rect 30172 25704 30732 25716
rect 31568 25750 31736 25762
rect 31568 25716 31574 25750
rect 31674 25716 31736 25750
rect 31960 25762 31972 26910
rect 32046 26726 33046 26830
rect 32046 25946 32156 26726
rect 32936 25946 33046 26726
rect 32046 25842 33046 25946
rect 33120 25762 33132 26910
rect 33356 27158 33368 28256
rect 34516 28256 34764 28306
rect 33442 28122 34442 28226
rect 33442 27342 33552 28122
rect 34332 27342 34442 28122
rect 33442 27238 34442 27342
rect 34516 27158 34528 28256
rect 33356 27146 33524 27158
rect 33356 27112 33418 27146
rect 33518 27112 33524 27146
rect 33356 27100 33524 27112
rect 34360 27146 34528 27158
rect 34360 27112 34366 27146
rect 34466 27112 34528 27146
rect 34360 27100 34528 27112
rect 33356 26968 33368 27100
rect 34516 26968 34528 27100
rect 33356 26956 33524 26968
rect 33356 26922 33418 26956
rect 33518 26922 33524 26956
rect 33356 26910 33524 26922
rect 34360 26956 34528 26968
rect 34360 26922 34366 26956
rect 34466 26922 34528 26956
rect 34360 26910 34528 26922
rect 31960 25750 32128 25762
rect 31960 25716 32022 25750
rect 32122 25716 32128 25750
rect 31568 25704 32128 25716
rect 32964 25750 33132 25762
rect 32964 25716 32970 25750
rect 33070 25716 33132 25750
rect 33356 25762 33368 26910
rect 33442 26726 34442 26830
rect 33442 25946 33552 26726
rect 34332 25946 34442 26726
rect 33442 25842 34442 25946
rect 34516 25762 34528 26910
rect 34752 27158 34764 28256
rect 35912 28256 36160 28306
rect 34838 28122 35838 28226
rect 34838 27342 34948 28122
rect 35728 27342 35838 28122
rect 34838 27238 35838 27342
rect 35912 27158 35924 28256
rect 34752 27146 34920 27158
rect 34752 27112 34814 27146
rect 34914 27112 34920 27146
rect 34752 27100 34920 27112
rect 35756 27146 35924 27158
rect 35756 27112 35762 27146
rect 35862 27112 35924 27146
rect 35756 27100 35924 27112
rect 34752 26968 34764 27100
rect 35912 26968 35924 27100
rect 34752 26956 34920 26968
rect 34752 26922 34814 26956
rect 34914 26922 34920 26956
rect 34752 26910 34920 26922
rect 35756 26956 35924 26968
rect 35756 26922 35762 26956
rect 35862 26922 35924 26956
rect 35756 26910 35924 26922
rect 33356 25750 33524 25762
rect 33356 25716 33418 25750
rect 33518 25716 33524 25750
rect 32964 25704 33524 25716
rect 34360 25750 34528 25762
rect 34360 25716 34366 25750
rect 34466 25716 34528 25750
rect 34752 25762 34764 26910
rect 34838 26726 35838 26830
rect 34838 25946 34948 26726
rect 35728 25946 35838 26726
rect 34838 25842 35838 25946
rect 35912 25762 35924 26910
rect 36148 27158 36160 28256
rect 37308 28256 37556 28306
rect 36234 28122 37234 28226
rect 36234 27342 36344 28122
rect 37124 27342 37234 28122
rect 36234 27238 37234 27342
rect 37308 27158 37320 28256
rect 36148 27146 36316 27158
rect 36148 27112 36210 27146
rect 36310 27112 36316 27146
rect 36148 27100 36316 27112
rect 37152 27146 37320 27158
rect 37152 27112 37158 27146
rect 37258 27112 37320 27146
rect 37152 27100 37320 27112
rect 36148 26968 36160 27100
rect 37308 26968 37320 27100
rect 36148 26956 36316 26968
rect 36148 26922 36210 26956
rect 36310 26922 36316 26956
rect 36148 26910 36316 26922
rect 37152 26956 37320 26968
rect 37152 26922 37158 26956
rect 37258 26922 37320 26956
rect 37152 26910 37320 26922
rect 34752 25750 34920 25762
rect 34752 25716 34814 25750
rect 34914 25716 34920 25750
rect 34360 25704 34920 25716
rect 35756 25750 35924 25762
rect 35756 25716 35762 25750
rect 35862 25716 35924 25750
rect 36148 25762 36160 26910
rect 36234 26726 37234 26830
rect 36234 25946 36344 26726
rect 37124 25946 37234 26726
rect 36234 25842 37234 25946
rect 37308 25762 37320 26910
rect 37544 27158 37556 28256
rect 38704 28256 38952 28306
rect 37630 28122 38630 28226
rect 37630 27342 37740 28122
rect 38520 27342 38630 28122
rect 37630 27238 38630 27342
rect 38704 27158 38716 28256
rect 37544 27146 37712 27158
rect 37544 27112 37606 27146
rect 37706 27112 37712 27146
rect 37544 27100 37712 27112
rect 38548 27146 38716 27158
rect 38548 27112 38554 27146
rect 38654 27112 38716 27146
rect 38548 27100 38716 27112
rect 37544 26968 37556 27100
rect 38704 26968 38716 27100
rect 37544 26956 37712 26968
rect 37544 26922 37606 26956
rect 37706 26922 37712 26956
rect 37544 26910 37712 26922
rect 38548 26956 38716 26968
rect 38548 26922 38554 26956
rect 38654 26922 38716 26956
rect 38548 26910 38716 26922
rect 36148 25750 36316 25762
rect 36148 25716 36210 25750
rect 36310 25716 36316 25750
rect 35756 25704 36316 25716
rect 37152 25750 37320 25762
rect 37152 25716 37158 25750
rect 37258 25716 37320 25750
rect 37544 25762 37556 26910
rect 37630 26726 38630 26830
rect 37630 25946 37740 26726
rect 38520 25946 38630 26726
rect 37630 25842 38630 25946
rect 38704 25762 38716 26910
rect 38940 27158 38952 28256
rect 40100 28256 40348 28306
rect 39026 28122 40026 28226
rect 39026 27342 39136 28122
rect 39916 27342 40026 28122
rect 39026 27238 40026 27342
rect 40100 27158 40112 28256
rect 38940 27146 39108 27158
rect 38940 27112 39002 27146
rect 39102 27112 39108 27146
rect 38940 27100 39108 27112
rect 39944 27146 40112 27158
rect 39944 27112 39950 27146
rect 40050 27112 40112 27146
rect 39944 27100 40112 27112
rect 38940 26968 38952 27100
rect 40100 26968 40112 27100
rect 38940 26956 39108 26968
rect 38940 26922 39002 26956
rect 39102 26922 39108 26956
rect 38940 26910 39108 26922
rect 39944 26956 40112 26968
rect 39944 26922 39950 26956
rect 40050 26922 40112 26956
rect 39944 26910 40112 26922
rect 37544 25750 37712 25762
rect 37544 25716 37606 25750
rect 37706 25716 37712 25750
rect 37152 25704 37712 25716
rect 38548 25750 38716 25762
rect 38548 25716 38554 25750
rect 38654 25716 38716 25750
rect 38940 25762 38952 26910
rect 39026 26726 40026 26830
rect 39026 25946 39136 26726
rect 39916 25946 40026 26726
rect 39026 25842 40026 25946
rect 40100 25762 40112 26910
rect 40336 27158 40348 28256
rect 41496 28256 41744 28306
rect 40422 28122 41422 28226
rect 40422 27342 40532 28122
rect 41312 27342 41422 28122
rect 40422 27238 41422 27342
rect 41496 27158 41508 28256
rect 40336 27146 40504 27158
rect 40336 27112 40398 27146
rect 40498 27112 40504 27146
rect 40336 27100 40504 27112
rect 41340 27146 41508 27158
rect 41340 27112 41346 27146
rect 41446 27112 41508 27146
rect 41340 27100 41508 27112
rect 40336 26968 40348 27100
rect 41496 26968 41508 27100
rect 40336 26956 40504 26968
rect 40336 26922 40398 26956
rect 40498 26922 40504 26956
rect 40336 26910 40504 26922
rect 41340 26956 41508 26968
rect 41340 26922 41346 26956
rect 41446 26922 41508 26956
rect 41340 26910 41508 26922
rect 38940 25750 39108 25762
rect 38940 25716 39002 25750
rect 39102 25716 39108 25750
rect 38548 25704 39108 25716
rect 39944 25750 40112 25762
rect 39944 25716 39950 25750
rect 40050 25716 40112 25750
rect 40336 25762 40348 26910
rect 40422 26726 41422 26830
rect 40422 25946 40532 26726
rect 41312 25946 41422 26726
rect 40422 25842 41422 25946
rect 41496 25762 41508 26910
rect 41732 27158 41744 28256
rect 42892 28256 43140 28306
rect 41818 28122 42818 28226
rect 41818 27342 41928 28122
rect 42708 27342 42818 28122
rect 41818 27238 42818 27342
rect 42892 27158 42904 28256
rect 41732 27146 41900 27158
rect 41732 27112 41794 27146
rect 41894 27112 41900 27146
rect 41732 27100 41900 27112
rect 42736 27146 42904 27158
rect 42736 27112 42742 27146
rect 42842 27112 42904 27146
rect 42736 27100 42904 27112
rect 41732 26968 41744 27100
rect 42892 26968 42904 27100
rect 41732 26956 41900 26968
rect 41732 26922 41794 26956
rect 41894 26922 41900 26956
rect 41732 26910 41900 26922
rect 42736 26956 42904 26968
rect 42736 26922 42742 26956
rect 42842 26922 42904 26956
rect 42736 26910 42904 26922
rect 40336 25750 40504 25762
rect 40336 25716 40398 25750
rect 40498 25716 40504 25750
rect 39944 25704 40504 25716
rect 41340 25750 41508 25762
rect 41340 25716 41346 25750
rect 41446 25716 41508 25750
rect 41732 25762 41744 26910
rect 41818 26726 42818 26830
rect 41818 25946 41928 26726
rect 42708 25946 42818 26726
rect 41818 25842 42818 25946
rect 42892 25762 42904 26910
rect 43128 27158 43140 28256
rect 44288 28256 44536 28306
rect 43214 28122 44214 28226
rect 43214 27342 43324 28122
rect 44104 27342 44214 28122
rect 43214 27238 44214 27342
rect 44288 27158 44300 28256
rect 43128 27146 43296 27158
rect 43128 27112 43190 27146
rect 43290 27112 43296 27146
rect 43128 27100 43296 27112
rect 44132 27146 44300 27158
rect 44132 27112 44138 27146
rect 44238 27112 44300 27146
rect 44132 27100 44300 27112
rect 43128 26968 43140 27100
rect 44288 26968 44300 27100
rect 43128 26956 43296 26968
rect 43128 26922 43190 26956
rect 43290 26922 43296 26956
rect 43128 26910 43296 26922
rect 44132 26956 44300 26968
rect 44132 26922 44138 26956
rect 44238 26922 44300 26956
rect 44132 26910 44300 26922
rect 41732 25750 41900 25762
rect 41732 25716 41794 25750
rect 41894 25716 41900 25750
rect 41340 25704 41900 25716
rect 42736 25750 42904 25762
rect 42736 25716 42742 25750
rect 42842 25716 42904 25750
rect 43128 25762 43140 26910
rect 43214 26726 44214 26830
rect 43214 25946 43324 26726
rect 44104 25946 44214 26726
rect 43214 25842 44214 25946
rect 44288 25762 44300 26910
rect 44524 27158 44536 28256
rect 45684 28256 45932 28306
rect 44610 28122 45610 28226
rect 44610 27342 44720 28122
rect 45500 27342 45610 28122
rect 44610 27238 45610 27342
rect 45684 27158 45696 28256
rect 44524 27146 44692 27158
rect 44524 27112 44586 27146
rect 44686 27112 44692 27146
rect 44524 27100 44692 27112
rect 45528 27146 45696 27158
rect 45528 27112 45534 27146
rect 45634 27112 45696 27146
rect 45528 27100 45696 27112
rect 44524 26968 44536 27100
rect 45684 26968 45696 27100
rect 44524 26956 44692 26968
rect 44524 26922 44586 26956
rect 44686 26922 44692 26956
rect 44524 26910 44692 26922
rect 45528 26956 45696 26968
rect 45528 26922 45534 26956
rect 45634 26922 45696 26956
rect 45528 26910 45696 26922
rect 43128 25750 43296 25762
rect 43128 25716 43190 25750
rect 43290 25716 43296 25750
rect 42736 25704 43296 25716
rect 44132 25750 44300 25762
rect 44132 25716 44138 25750
rect 44238 25716 44300 25750
rect 44524 25762 44536 26910
rect 44610 26726 45610 26830
rect 44610 25946 44720 26726
rect 45500 25946 45610 26726
rect 44610 25842 45610 25946
rect 45684 25762 45696 26910
rect 45920 27158 45932 28256
rect 47080 28256 47328 28306
rect 46006 28122 47006 28226
rect 46006 27342 46116 28122
rect 46896 27342 47006 28122
rect 46006 27238 47006 27342
rect 47080 27158 47092 28256
rect 45920 27146 46088 27158
rect 45920 27112 45982 27146
rect 46082 27112 46088 27146
rect 45920 27100 46088 27112
rect 46924 27146 47092 27158
rect 46924 27112 46930 27146
rect 47030 27112 47092 27146
rect 46924 27100 47092 27112
rect 45920 26968 45932 27100
rect 47080 26968 47092 27100
rect 45920 26956 46088 26968
rect 45920 26922 45982 26956
rect 46082 26922 46088 26956
rect 45920 26910 46088 26922
rect 46924 26956 47092 26968
rect 46924 26922 46930 26956
rect 47030 26922 47092 26956
rect 46924 26910 47092 26922
rect 44524 25750 44692 25762
rect 44524 25716 44586 25750
rect 44686 25716 44692 25750
rect 44132 25704 44692 25716
rect 45528 25750 45696 25762
rect 45528 25716 45534 25750
rect 45634 25716 45696 25750
rect 45920 25762 45932 26910
rect 46006 26726 47006 26830
rect 46006 25946 46116 26726
rect 46896 25946 47006 26726
rect 46006 25842 47006 25946
rect 47080 25762 47092 26910
rect 47316 27158 47328 28256
rect 48476 28256 48724 28306
rect 47402 28122 48402 28226
rect 47402 27342 47512 28122
rect 48292 27342 48402 28122
rect 47402 27238 48402 27342
rect 48476 27158 48488 28256
rect 47316 27146 47484 27158
rect 47316 27112 47378 27146
rect 47478 27112 47484 27146
rect 47316 27100 47484 27112
rect 48320 27146 48488 27158
rect 48320 27112 48326 27146
rect 48426 27112 48488 27146
rect 48320 27100 48488 27112
rect 47316 26968 47328 27100
rect 48476 26968 48488 27100
rect 47316 26956 47484 26968
rect 47316 26922 47378 26956
rect 47478 26922 47484 26956
rect 47316 26910 47484 26922
rect 48320 26956 48488 26968
rect 48320 26922 48326 26956
rect 48426 26922 48488 26956
rect 48320 26910 48488 26922
rect 45920 25750 46088 25762
rect 45920 25716 45982 25750
rect 46082 25716 46088 25750
rect 45528 25704 46088 25716
rect 46924 25750 47092 25762
rect 46924 25716 46930 25750
rect 47030 25716 47092 25750
rect 47316 25762 47328 26910
rect 47402 26726 48402 26830
rect 47402 25946 47512 26726
rect 48292 25946 48402 26726
rect 47402 25842 48402 25946
rect 48476 25762 48488 26910
rect 48712 27158 48724 28256
rect 49872 28256 50120 28306
rect 48798 28122 49798 28226
rect 48798 27342 48908 28122
rect 49688 27342 49798 28122
rect 48798 27238 49798 27342
rect 49872 27158 49884 28256
rect 48712 27146 48880 27158
rect 48712 27112 48774 27146
rect 48874 27112 48880 27146
rect 48712 27100 48880 27112
rect 49716 27146 49884 27158
rect 49716 27112 49722 27146
rect 49822 27112 49884 27146
rect 49716 27100 49884 27112
rect 48712 26968 48724 27100
rect 49872 26968 49884 27100
rect 48712 26956 48880 26968
rect 48712 26922 48774 26956
rect 48874 26922 48880 26956
rect 48712 26910 48880 26922
rect 49716 26956 49884 26968
rect 49716 26922 49722 26956
rect 49822 26922 49884 26956
rect 49716 26910 49884 26922
rect 47316 25750 47484 25762
rect 47316 25716 47378 25750
rect 47478 25716 47484 25750
rect 46924 25704 47484 25716
rect 48320 25750 48488 25762
rect 48320 25716 48326 25750
rect 48426 25716 48488 25750
rect 48712 25762 48724 26910
rect 48798 26726 49798 26830
rect 48798 25946 48908 26726
rect 49688 25946 49798 26726
rect 48798 25842 49798 25946
rect 49872 25762 49884 26910
rect 50108 27158 50120 28256
rect 51268 28256 51392 28306
rect 50194 28122 51194 28226
rect 50194 27342 50304 28122
rect 51084 27342 51194 28122
rect 50194 27238 51194 27342
rect 51268 27208 51280 28256
rect 51314 27208 51392 28256
rect 51268 27158 51392 27208
rect 50108 27146 50276 27158
rect 50108 27112 50170 27146
rect 50270 27112 50276 27146
rect 50108 27100 50276 27112
rect 51112 27146 51392 27158
rect 51112 27112 51118 27146
rect 51218 27112 51392 27146
rect 51112 27100 51392 27112
rect 50108 26968 50120 27100
rect 51268 26968 51392 27100
rect 50108 26956 50276 26968
rect 50108 26922 50170 26956
rect 50270 26922 50276 26956
rect 50108 26910 50276 26922
rect 51112 26956 51392 26968
rect 51112 26922 51118 26956
rect 51218 26922 51392 26956
rect 51112 26910 51392 26922
rect 48712 25750 48880 25762
rect 48712 25716 48774 25750
rect 48874 25716 48880 25750
rect 48320 25704 48880 25716
rect 49716 25750 49884 25762
rect 49716 25716 49722 25750
rect 49822 25716 49884 25750
rect 50108 25762 50120 26910
rect 51268 26860 51392 26910
rect 50194 26726 51194 26830
rect 50194 25946 50304 26726
rect 51084 25946 51194 26726
rect 50194 25842 51194 25946
rect 51268 25812 51280 26860
rect 51314 25812 51392 26860
rect 51268 25762 51392 25812
rect 50108 25750 50276 25762
rect 50108 25716 50170 25750
rect 50270 25716 50276 25750
rect 49716 25704 50276 25716
rect 51112 25750 51392 25762
rect 51112 25716 51118 25750
rect 51218 25716 51392 25750
rect 51112 25704 51392 25716
rect 9368 25552 9426 25602
rect 51478 25602 51490 28466
rect 51524 25846 51536 28466
rect 51524 25646 70826 25846
rect 51524 25602 51536 25646
rect 51478 25552 51536 25602
rect 9368 25540 51536 25552
rect 9368 25506 9476 25540
rect 51428 25506 51536 25540
rect 9368 25494 51536 25506
rect 3928 24928 4298 24978
rect -1780 24918 4298 24928
rect -1780 24690 -1696 24918
rect -1368 24916 -300 24918
rect -1368 24882 -1358 24916
rect -310 24882 -300 24916
rect -1368 24690 -300 24882
rect 28 24916 1096 24918
rect 28 24882 38 24916
rect 1086 24882 1096 24916
rect 28 24690 1096 24882
rect 1424 24916 2492 24918
rect 1424 24882 1434 24916
rect 2482 24882 2492 24916
rect 1424 24690 2492 24882
rect 2820 24916 3888 24918
rect 2820 24882 2830 24916
rect 3878 24882 3888 24916
rect 2820 24690 3888 24882
rect 4216 24690 4298 24918
rect -18962 24458 -3762 24646
rect -1780 24558 4298 24690
rect -1780 24556 4280 24558
rect -18962 23250 -18362 24458
rect -17410 24278 -17216 24284
rect -17792 24054 -17584 24062
rect -17792 23654 -17786 24054
rect -17590 23654 -17584 24054
rect -17792 23648 -17584 23654
rect -17410 23436 -17404 24278
rect -17222 23436 -17216 24278
rect -17410 23430 -17216 23436
rect -17184 23250 -16786 24458
rect -16004 24278 -15810 24284
rect -16386 24054 -16178 24062
rect -16386 23654 -16380 24054
rect -16184 23654 -16178 24054
rect -16386 23648 -16178 23654
rect -16004 23436 -15998 24278
rect -15816 23436 -15810 24278
rect -16004 23430 -15810 23436
rect -15778 23250 -15380 24458
rect -14598 24278 -14404 24284
rect -14980 24054 -14772 24062
rect -14980 23654 -14974 24054
rect -14778 23654 -14772 24054
rect -14980 23648 -14772 23654
rect -14598 23436 -14592 24278
rect -14410 23436 -14404 24278
rect -14598 23430 -14404 23436
rect -14372 23250 -13974 24458
rect -13192 24278 -12998 24284
rect -13574 24054 -13366 24062
rect -13574 23654 -13568 24054
rect -13372 23654 -13366 24054
rect -13574 23648 -13366 23654
rect -13192 23436 -13186 24278
rect -13004 23436 -12998 24278
rect -13192 23430 -12998 23436
rect -12966 23250 -12568 24458
rect -11786 24278 -11592 24284
rect -12168 24054 -11960 24062
rect -12168 23654 -12162 24054
rect -11966 23654 -11960 24054
rect -12168 23648 -11960 23654
rect -11786 23436 -11780 24278
rect -11598 23436 -11592 24278
rect -11786 23430 -11592 23436
rect -11560 23250 -11162 24458
rect -10380 24278 -10186 24284
rect -10762 24054 -10554 24062
rect -10762 23654 -10756 24054
rect -10560 23654 -10554 24054
rect -10762 23648 -10554 23654
rect -10380 23436 -10374 24278
rect -10192 23436 -10186 24278
rect -10380 23430 -10186 23436
rect -10154 23250 -9756 24458
rect -8974 24278 -8780 24284
rect -9356 24054 -9148 24062
rect -9356 23654 -9350 24054
rect -9154 23654 -9148 24054
rect -9356 23648 -9148 23654
rect -8974 23436 -8968 24278
rect -8786 23436 -8780 24278
rect -8974 23430 -8780 23436
rect -8748 23250 -8350 24458
rect -7568 24278 -7374 24284
rect -7950 24054 -7742 24062
rect -7950 23654 -7944 24054
rect -7748 23654 -7742 24054
rect -7950 23648 -7742 23654
rect -7568 23436 -7562 24278
rect -7380 23436 -7374 24278
rect -7568 23430 -7374 23436
rect -7342 23250 -6944 24458
rect -6162 24278 -5968 24284
rect -6544 24054 -6336 24062
rect -6544 23654 -6538 24054
rect -6342 23654 -6336 24054
rect -6544 23648 -6336 23654
rect -6162 23436 -6156 24278
rect -5974 23436 -5968 24278
rect -6162 23430 -5968 23436
rect -5936 23250 -5538 24458
rect -4362 24446 -3762 24458
rect -4362 24438 3628 24446
rect -4756 24278 -4562 24284
rect -5138 24054 -4930 24062
rect -5138 23654 -5132 24054
rect -4936 23654 -4930 24054
rect -5138 23648 -4930 23654
rect -4756 23436 -4750 24278
rect -4568 23436 -4562 24278
rect -4756 23430 -4562 23436
rect -4362 23856 -1228 24438
rect 3618 23856 3628 24438
rect -4362 23846 3628 23856
rect 3698 24414 4098 24432
rect 3698 24054 3718 24414
rect 4078 24054 4098 24414
rect -4362 23646 -3762 23846
rect -732 23646 -132 23846
rect -4362 23250 -132 23646
rect -18962 23046 -132 23250
rect -18962 22852 -3762 23046
rect -18962 21644 -18362 22852
rect -17410 22672 -17216 22678
rect -17792 22448 -17584 22456
rect -17792 22048 -17786 22448
rect -17590 22048 -17584 22448
rect -17792 22042 -17584 22048
rect -17410 21830 -17404 22672
rect -17222 21830 -17216 22672
rect -17410 21824 -17216 21830
rect -17184 21644 -16786 22852
rect -16004 22672 -15810 22678
rect -16386 22448 -16178 22456
rect -16386 22048 -16380 22448
rect -16184 22048 -16178 22448
rect -16386 22042 -16178 22048
rect -16004 21830 -15998 22672
rect -15816 21830 -15810 22672
rect -16004 21824 -15810 21830
rect -15778 21644 -15380 22852
rect -14598 22672 -14404 22678
rect -14980 22448 -14772 22456
rect -14980 22048 -14974 22448
rect -14778 22048 -14772 22448
rect -14980 22042 -14772 22048
rect -14598 21830 -14592 22672
rect -14410 21830 -14404 22672
rect -14598 21824 -14404 21830
rect -14372 21644 -13974 22852
rect -13192 22672 -12998 22678
rect -13574 22448 -13366 22456
rect -13574 22048 -13568 22448
rect -13372 22048 -13366 22448
rect -13574 22042 -13366 22048
rect -13192 21830 -13186 22672
rect -13004 21830 -12998 22672
rect -13192 21824 -12998 21830
rect -12966 21644 -12568 22852
rect -11786 22672 -11592 22678
rect -12168 22448 -11960 22456
rect -12168 22048 -12162 22448
rect -11966 22048 -11960 22448
rect -12168 22042 -11960 22048
rect -11786 21830 -11780 22672
rect -11598 21830 -11592 22672
rect -11786 21824 -11592 21830
rect -11560 21644 -11162 22852
rect -10380 22672 -10186 22678
rect -10762 22448 -10554 22456
rect -10762 22048 -10756 22448
rect -10560 22048 -10554 22448
rect -10762 22042 -10554 22048
rect -10380 21830 -10374 22672
rect -10192 21830 -10186 22672
rect -10380 21824 -10186 21830
rect -10154 21644 -9756 22852
rect -8974 22672 -8780 22678
rect -9356 22448 -9148 22456
rect -9356 22048 -9350 22448
rect -9154 22048 -9148 22448
rect -9356 22042 -9148 22048
rect -8974 21830 -8968 22672
rect -8786 21830 -8780 22672
rect -8974 21824 -8780 21830
rect -8748 21644 -8350 22852
rect -7568 22672 -7374 22678
rect -7950 22448 -7742 22456
rect -7950 22048 -7944 22448
rect -7748 22048 -7742 22448
rect -7950 22042 -7742 22048
rect -7568 21830 -7562 22672
rect -7380 21830 -7374 22672
rect -7568 21824 -7374 21830
rect -7342 21644 -6944 22852
rect -6162 22672 -5968 22678
rect -6544 22448 -6336 22456
rect -6544 22048 -6538 22448
rect -6342 22048 -6336 22448
rect -6544 22042 -6336 22048
rect -6162 21830 -6156 22672
rect -5974 21830 -5968 22672
rect -6162 21824 -5968 21830
rect -5936 21644 -5538 22852
rect -4362 22846 -3762 22852
rect 68 22846 668 23846
rect -4756 22672 -4562 22678
rect -5138 22448 -4930 22456
rect -5138 22048 -5132 22448
rect -4936 22048 -4930 22448
rect -5138 22042 -4930 22048
rect -4756 21830 -4750 22672
rect -4568 21830 -4562 22672
rect -4756 21824 -4562 21830
rect -4362 22246 668 22846
rect -4362 22046 -3762 22246
rect 868 22046 1468 23846
rect -4362 21644 1468 22046
rect -18962 21446 1468 21644
rect -18962 21246 -3762 21446
rect 1668 21246 2268 23846
rect -18962 20038 -18362 21246
rect -17410 21066 -17216 21072
rect -17792 20842 -17584 20850
rect -17792 20442 -17786 20842
rect -17590 20442 -17584 20842
rect -17792 20436 -17584 20442
rect -17410 20224 -17404 21066
rect -17222 20224 -17216 21066
rect -17410 20218 -17216 20224
rect -17184 20038 -16786 21246
rect -16004 21066 -15810 21072
rect -16386 20842 -16178 20850
rect -16386 20442 -16380 20842
rect -16184 20442 -16178 20842
rect -16386 20436 -16178 20442
rect -16004 20224 -15998 21066
rect -15816 20224 -15810 21066
rect -16004 20218 -15810 20224
rect -15778 20038 -15380 21246
rect -14598 21066 -14404 21072
rect -14980 20842 -14772 20850
rect -14980 20442 -14974 20842
rect -14778 20442 -14772 20842
rect -14980 20436 -14772 20442
rect -14598 20224 -14592 21066
rect -14410 20224 -14404 21066
rect -14598 20218 -14404 20224
rect -14372 20038 -13974 21246
rect -13192 21066 -12998 21072
rect -13574 20842 -13366 20850
rect -13574 20442 -13568 20842
rect -13372 20442 -13366 20842
rect -13574 20436 -13366 20442
rect -13192 20224 -13186 21066
rect -13004 20224 -12998 21066
rect -13192 20218 -12998 20224
rect -12966 20038 -12568 21246
rect -11786 21066 -11592 21072
rect -12168 20842 -11960 20850
rect -12168 20442 -12162 20842
rect -11966 20442 -11960 20842
rect -12168 20436 -11960 20442
rect -11786 20224 -11780 21066
rect -11598 20224 -11592 21066
rect -11786 20218 -11592 20224
rect -11560 20038 -11162 21246
rect -10380 21066 -10186 21072
rect -10762 20842 -10554 20850
rect -10762 20442 -10756 20842
rect -10560 20442 -10554 20842
rect -10762 20436 -10554 20442
rect -10380 20224 -10374 21066
rect -10192 20224 -10186 21066
rect -10380 20218 -10186 20224
rect -10154 20038 -9756 21246
rect -8974 21066 -8780 21072
rect -9356 20842 -9148 20850
rect -9356 20442 -9350 20842
rect -9154 20442 -9148 20842
rect -9356 20436 -9148 20442
rect -8974 20224 -8968 21066
rect -8786 20224 -8780 21066
rect -8974 20218 -8780 20224
rect -8748 20038 -8350 21246
rect -7568 21066 -7374 21072
rect -7950 20842 -7742 20850
rect -7950 20442 -7944 20842
rect -7748 20442 -7742 20842
rect -7950 20436 -7742 20442
rect -7568 20224 -7562 21066
rect -7380 20224 -7374 21066
rect -7568 20218 -7374 20224
rect -7342 20038 -6944 21246
rect -6162 21066 -5968 21072
rect -6544 20842 -6336 20850
rect -6544 20442 -6538 20842
rect -6342 20442 -6336 20842
rect -6544 20436 -6336 20442
rect -6162 20224 -6156 21066
rect -5974 20224 -5968 21066
rect -6162 20218 -5968 20224
rect -5936 20038 -5538 21246
rect -4756 21066 -4562 21072
rect -5138 20842 -4930 20850
rect -5138 20442 -5132 20842
rect -4936 20442 -4930 20842
rect -5138 20436 -4930 20442
rect -4756 20224 -4750 21066
rect -4568 20224 -4562 21066
rect -4756 20218 -4562 20224
rect -4362 20646 2268 21246
rect -4362 20446 -3762 20646
rect 2468 20446 3068 23846
rect 3698 23344 4098 24054
rect 3690 23336 4106 23344
rect 3690 22936 3698 23336
rect 4098 22936 4106 23336
rect 3690 22928 4106 22936
rect -4362 20038 3068 20446
rect -18962 19846 3068 20038
rect -18962 19640 -3762 19846
rect -18962 18432 -18362 19640
rect -17410 19460 -17216 19466
rect -17792 19236 -17584 19244
rect -17792 18836 -17786 19236
rect -17590 18836 -17584 19236
rect -17792 18830 -17584 18836
rect -17410 18618 -17404 19460
rect -17222 18618 -17216 19460
rect -17410 18612 -17216 18618
rect -17184 18432 -16786 19640
rect -16004 19460 -15810 19466
rect -16386 19236 -16178 19244
rect -16386 18836 -16380 19236
rect -16184 18836 -16178 19236
rect -16386 18830 -16178 18836
rect -16004 18618 -15998 19460
rect -15816 18618 -15810 19460
rect -16004 18612 -15810 18618
rect -15778 18432 -15380 19640
rect -14598 19460 -14404 19466
rect -14980 19236 -14772 19244
rect -14980 18836 -14974 19236
rect -14778 18836 -14772 19236
rect -14980 18830 -14772 18836
rect -14598 18618 -14592 19460
rect -14410 18618 -14404 19460
rect -14598 18612 -14404 18618
rect -14372 18432 -13974 19640
rect -13192 19460 -12998 19466
rect -13574 19236 -13366 19244
rect -13574 18836 -13568 19236
rect -13372 18836 -13366 19236
rect -13574 18830 -13366 18836
rect -13192 18618 -13186 19460
rect -13004 18618 -12998 19460
rect -13192 18612 -12998 18618
rect -12966 18432 -12568 19640
rect -11786 19460 -11592 19466
rect -12168 19236 -11960 19244
rect -12168 18836 -12162 19236
rect -11966 18836 -11960 19236
rect -12168 18830 -11960 18836
rect -11786 18618 -11780 19460
rect -11598 18618 -11592 19460
rect -11786 18612 -11592 18618
rect -11560 18432 -11162 19640
rect -10380 19460 -10186 19466
rect -10762 19236 -10554 19244
rect -10762 18836 -10756 19236
rect -10560 18836 -10554 19236
rect -10762 18830 -10554 18836
rect -10380 18618 -10374 19460
rect -10192 18618 -10186 19460
rect -10380 18612 -10186 18618
rect -10154 18432 -9756 19640
rect -8974 19460 -8780 19466
rect -9356 19236 -9148 19244
rect -9356 18836 -9350 19236
rect -9154 18836 -9148 19236
rect -9356 18830 -9148 18836
rect -8974 18618 -8968 19460
rect -8786 18618 -8780 19460
rect -8974 18612 -8780 18618
rect -8748 18432 -8350 19640
rect -7568 19460 -7374 19466
rect -7950 19236 -7742 19244
rect -7950 18836 -7944 19236
rect -7748 18836 -7742 19236
rect -7950 18830 -7742 18836
rect -7568 18618 -7562 19460
rect -7380 18618 -7374 19460
rect -7568 18612 -7374 18618
rect -7342 18432 -6944 19640
rect -6162 19460 -5968 19466
rect -6544 19236 -6336 19244
rect -6544 18836 -6538 19236
rect -6342 18836 -6336 19236
rect -6544 18830 -6336 18836
rect -6162 18618 -6156 19460
rect -5974 18618 -5968 19460
rect -6162 18612 -5968 18618
rect -5936 18432 -5538 19640
rect -4756 19460 -4562 19466
rect -5138 19236 -4930 19244
rect -5138 18836 -5132 19236
rect -4936 18836 -4930 19236
rect -5138 18830 -4930 18836
rect -4756 18618 -4750 19460
rect -4568 18618 -4562 19460
rect -4756 18612 -4562 18618
rect -4362 18432 -3762 19640
rect -2980 19040 -2560 19048
rect -2980 18640 -2968 19040
rect -2568 18640 -2560 19040
rect -2980 18630 -2560 18640
rect -18962 18034 -3762 18432
rect -18962 16826 -18362 18034
rect -17410 17854 -17216 17860
rect -17792 17630 -17584 17638
rect -17792 17230 -17786 17630
rect -17590 17230 -17584 17630
rect -17792 17224 -17584 17230
rect -17410 17012 -17404 17854
rect -17222 17012 -17216 17854
rect -17410 17006 -17216 17012
rect -17184 16826 -16786 18034
rect -16004 17854 -15810 17860
rect -16386 17630 -16178 17638
rect -16386 17230 -16380 17630
rect -16184 17230 -16178 17630
rect -16386 17224 -16178 17230
rect -16004 17012 -15998 17854
rect -15816 17012 -15810 17854
rect -16004 17006 -15810 17012
rect -15778 16826 -15380 18034
rect -14598 17854 -14404 17860
rect -14980 17630 -14772 17638
rect -14980 17230 -14974 17630
rect -14778 17230 -14772 17630
rect -14980 17224 -14772 17230
rect -14598 17012 -14592 17854
rect -14410 17012 -14404 17854
rect -14598 17006 -14404 17012
rect -14372 16826 -13974 18034
rect -13192 17854 -12998 17860
rect -13574 17630 -13366 17638
rect -13574 17230 -13568 17630
rect -13372 17230 -13366 17630
rect -13574 17224 -13366 17230
rect -13192 17012 -13186 17854
rect -13004 17012 -12998 17854
rect -13192 17006 -12998 17012
rect -12966 16826 -12568 18034
rect -11786 17854 -11592 17860
rect -12168 17630 -11960 17638
rect -12168 17230 -12162 17630
rect -11966 17230 -11960 17630
rect -12168 17224 -11960 17230
rect -11786 17012 -11780 17854
rect -11598 17012 -11592 17854
rect -11786 17006 -11592 17012
rect -11560 16826 -11162 18034
rect -10380 17854 -10186 17860
rect -10762 17630 -10554 17638
rect -10762 17230 -10756 17630
rect -10560 17230 -10554 17630
rect -10762 17224 -10554 17230
rect -10380 17012 -10374 17854
rect -10192 17012 -10186 17854
rect -10380 17006 -10186 17012
rect -10154 16826 -9756 18034
rect -8974 17854 -8780 17860
rect -9356 17630 -9148 17638
rect -9356 17230 -9350 17630
rect -9154 17230 -9148 17630
rect -9356 17224 -9148 17230
rect -8974 17012 -8968 17854
rect -8786 17012 -8780 17854
rect -8974 17006 -8780 17012
rect -8748 16826 -8350 18034
rect -7568 17854 -7374 17860
rect -7950 17630 -7742 17638
rect -7950 17230 -7944 17630
rect -7748 17230 -7742 17630
rect -7950 17224 -7742 17230
rect -7568 17012 -7562 17854
rect -7380 17012 -7374 17854
rect -7568 17006 -7374 17012
rect -7342 16826 -6944 18034
rect -6162 17854 -5968 17860
rect -6544 17630 -6336 17638
rect -6544 17230 -6538 17630
rect -6342 17230 -6336 17630
rect -6544 17224 -6336 17230
rect -6162 17012 -6156 17854
rect -5974 17012 -5968 17854
rect -6162 17006 -5968 17012
rect -5936 16826 -5538 18034
rect -4756 17854 -4562 17860
rect -5138 17630 -4930 17638
rect -5138 17230 -5132 17630
rect -4936 17230 -4930 17630
rect -5138 17224 -4930 17230
rect -4756 17012 -4750 17854
rect -4568 17012 -4562 17854
rect -4756 17006 -4562 17012
rect -4362 16826 -3762 18034
rect -18962 16428 -3762 16826
rect -18962 15220 -18362 16428
rect -17410 16248 -17216 16254
rect -17792 16024 -17584 16032
rect -17792 15624 -17786 16024
rect -17590 15624 -17584 16024
rect -17792 15618 -17584 15624
rect -17410 15406 -17404 16248
rect -17222 15406 -17216 16248
rect -17410 15400 -17216 15406
rect -17184 15220 -16786 16428
rect -16004 16248 -15810 16254
rect -16386 16024 -16178 16032
rect -16386 15624 -16380 16024
rect -16184 15624 -16178 16024
rect -16386 15618 -16178 15624
rect -16004 15406 -15998 16248
rect -15816 15406 -15810 16248
rect -16004 15400 -15810 15406
rect -15778 15220 -15380 16428
rect -14598 16248 -14404 16254
rect -14980 16024 -14772 16032
rect -14980 15624 -14974 16024
rect -14778 15624 -14772 16024
rect -14980 15618 -14772 15624
rect -14598 15406 -14592 16248
rect -14410 15406 -14404 16248
rect -14598 15400 -14404 15406
rect -14372 15220 -13974 16428
rect -13192 16248 -12998 16254
rect -13574 16024 -13366 16032
rect -13574 15624 -13568 16024
rect -13372 15624 -13366 16024
rect -13574 15618 -13366 15624
rect -13192 15406 -13186 16248
rect -13004 15406 -12998 16248
rect -13192 15400 -12998 15406
rect -12966 15220 -12568 16428
rect -11786 16248 -11592 16254
rect -12168 16024 -11960 16032
rect -12168 15624 -12162 16024
rect -11966 15624 -11960 16024
rect -12168 15618 -11960 15624
rect -11786 15406 -11780 16248
rect -11598 15406 -11592 16248
rect -11786 15400 -11592 15406
rect -11560 15220 -11162 16428
rect -10380 16248 -10186 16254
rect -10762 16024 -10554 16032
rect -10762 15624 -10756 16024
rect -10560 15624 -10554 16024
rect -10762 15618 -10554 15624
rect -10380 15406 -10374 16248
rect -10192 15406 -10186 16248
rect -10380 15400 -10186 15406
rect -10154 15220 -9756 16428
rect -8974 16248 -8780 16254
rect -9356 16024 -9148 16032
rect -9356 15624 -9350 16024
rect -9154 15624 -9148 16024
rect -9356 15618 -9148 15624
rect -8974 15406 -8968 16248
rect -8786 15406 -8780 16248
rect -8974 15400 -8780 15406
rect -8748 15220 -8350 16428
rect -7568 16248 -7374 16254
rect -7950 16024 -7742 16032
rect -7950 15624 -7944 16024
rect -7748 15624 -7742 16024
rect -7950 15618 -7742 15624
rect -7568 15406 -7562 16248
rect -7380 15406 -7374 16248
rect -7568 15400 -7374 15406
rect -7342 15220 -6944 16428
rect -6162 16248 -5968 16254
rect -6544 16024 -6336 16032
rect -6544 15624 -6538 16024
rect -6342 15624 -6336 16024
rect -6544 15618 -6336 15624
rect -6162 15406 -6156 16248
rect -5974 15406 -5968 16248
rect -6162 15400 -5968 15406
rect -5936 15220 -5538 16428
rect -4756 16248 -4562 16254
rect -5138 16024 -4930 16032
rect -5138 15624 -5132 16024
rect -4936 15624 -4930 16024
rect -5138 15618 -4930 15624
rect -4756 15406 -4750 16248
rect -4568 15406 -4562 16248
rect -4756 15400 -4562 15406
rect -4362 15220 -3762 16428
rect -18962 14822 -3762 15220
rect -18962 13504 -18362 14822
rect -17410 14642 -17216 14648
rect -17792 14418 -17584 14426
rect -17792 14018 -17786 14418
rect -17590 14018 -17584 14418
rect -17792 14012 -17584 14018
rect -17410 13800 -17404 14642
rect -17222 13800 -17216 14642
rect -17410 13794 -17216 13800
rect -17184 13504 -16786 14822
rect -16004 14642 -15810 14648
rect -16386 14418 -16178 14426
rect -16386 14018 -16380 14418
rect -16184 14018 -16178 14418
rect -16386 14012 -16178 14018
rect -16004 13800 -15998 14642
rect -15816 13800 -15810 14642
rect -16004 13794 -15810 13800
rect -15778 13504 -15380 14822
rect -14598 14642 -14404 14648
rect -14980 14418 -14772 14426
rect -14980 14018 -14974 14418
rect -14778 14018 -14772 14418
rect -14980 14012 -14772 14018
rect -14598 13800 -14592 14642
rect -14410 13800 -14404 14642
rect -14598 13794 -14404 13800
rect -14372 13504 -13974 14822
rect -13192 14642 -12998 14648
rect -13574 14418 -13366 14426
rect -13574 14018 -13568 14418
rect -13372 14018 -13366 14418
rect -13574 14012 -13366 14018
rect -13192 13800 -13186 14642
rect -13004 13800 -12998 14642
rect -13192 13794 -12998 13800
rect -12966 13504 -12568 14822
rect -11786 14642 -11592 14648
rect -12168 14418 -11960 14426
rect -12168 14018 -12162 14418
rect -11966 14018 -11960 14418
rect -12168 14012 -11960 14018
rect -11786 13800 -11780 14642
rect -11598 13800 -11592 14642
rect -11786 13794 -11592 13800
rect -11560 13504 -11162 14822
rect -10380 14642 -10186 14648
rect -10762 14418 -10554 14426
rect -10762 14018 -10756 14418
rect -10560 14018 -10554 14418
rect -10762 14012 -10554 14018
rect -10380 13800 -10374 14642
rect -10192 13800 -10186 14642
rect -10380 13794 -10186 13800
rect -10154 13504 -9756 14822
rect -8974 14642 -8780 14648
rect -9356 14418 -9148 14426
rect -9356 14018 -9350 14418
rect -9154 14018 -9148 14418
rect -9356 14012 -9148 14018
rect -8974 13800 -8968 14642
rect -8786 13800 -8780 14642
rect -8974 13794 -8780 13800
rect -8748 13504 -8350 14822
rect -7568 14642 -7374 14648
rect -7950 14418 -7742 14426
rect -7950 14018 -7944 14418
rect -7748 14018 -7742 14418
rect -7950 14012 -7742 14018
rect -7568 13800 -7562 14642
rect -7380 13800 -7374 14642
rect -7568 13794 -7374 13800
rect -7342 13504 -6944 14822
rect -6162 14642 -5968 14648
rect -6544 14418 -6336 14426
rect -6544 14018 -6538 14418
rect -6342 14018 -6336 14418
rect -6544 14012 -6336 14018
rect -6162 13800 -6156 14642
rect -5974 13800 -5968 14642
rect -6162 13794 -5968 13800
rect -5936 13504 -5538 14822
rect -4756 14642 -4562 14648
rect -5138 14418 -4930 14426
rect -5138 14018 -5132 14418
rect -4936 14018 -4930 14418
rect -5138 14012 -4930 14018
rect -4756 13800 -4750 14642
rect -4568 13800 -4562 14642
rect -4756 13794 -4562 13800
rect -4362 13504 -3762 14822
rect -18962 12904 -3762 13504
rect 526 13428 616 13434
rect 842 13428 932 13434
rect 1158 13428 1248 13434
rect 1474 13428 1564 13434
rect 1790 13428 1880 13438
rect 2106 13428 2196 13438
rect 2422 13428 2512 13434
rect 2738 13428 2828 13434
rect 3054 13428 3144 13434
rect 3370 13428 3460 13434
rect 250 13426 3740 13428
rect 250 13412 538 13426
rect 3448 13412 3740 13426
rect 250 13378 360 13412
rect 3630 13378 3740 13412
rect 250 13370 538 13378
rect 3448 13370 3740 13378
rect 250 13362 3740 13370
rect 250 13316 314 13362
rect 526 13358 616 13362
rect 842 13358 932 13362
rect 1158 13358 1248 13362
rect 1474 13358 1564 13362
rect 1790 13358 1880 13362
rect 2106 13358 2196 13362
rect 2422 13358 2512 13362
rect 2738 13358 2828 13362
rect 3054 13358 3144 13362
rect 3370 13358 3460 13362
rect 250 12074 264 13316
rect 298 12074 314 13316
rect 3676 13316 3740 13362
rect 378 13242 3598 13300
rect 380 13234 3598 13242
rect 380 12970 438 13234
rect 540 13202 606 13206
rect 540 13004 546 13202
rect 600 13004 606 13202
rect 540 12998 606 13004
rect 708 12970 754 13234
rect 856 13202 922 13206
rect 856 13004 862 13202
rect 916 13004 922 13202
rect 856 12998 922 13004
rect 1024 12970 1070 13234
rect 1172 13202 1238 13206
rect 1172 13004 1178 13202
rect 1232 13004 1238 13202
rect 1172 12998 1238 13004
rect 1340 12970 1386 13234
rect 1488 13202 1554 13206
rect 1488 13004 1494 13202
rect 1548 13004 1554 13202
rect 1488 12998 1554 13004
rect 1656 12970 1702 13234
rect 1804 13202 1870 13206
rect 1804 13004 1810 13202
rect 1864 13004 1870 13202
rect 1804 12998 1870 13004
rect 1972 12970 2018 13234
rect 2120 13202 2186 13206
rect 2120 13004 2126 13202
rect 2180 13004 2186 13202
rect 2120 12998 2186 13004
rect 2288 12970 2334 13234
rect 2436 13202 2502 13206
rect 2436 13004 2442 13202
rect 2496 13004 2502 13202
rect 2436 12998 2502 13004
rect 2604 12970 2650 13234
rect 2752 13202 2818 13206
rect 2752 13004 2758 13202
rect 2812 13004 2818 13202
rect 2752 12998 2818 13004
rect 2920 12970 2966 13234
rect 3068 13202 3134 13206
rect 3068 13004 3074 13202
rect 3128 13004 3134 13202
rect 3068 12998 3134 13004
rect 3236 12970 3282 13234
rect 3384 13202 3450 13206
rect 3384 13004 3390 13202
rect 3444 13004 3450 13202
rect 3384 12998 3450 13004
rect 3550 12970 3598 13234
rect 380 12968 3598 12970
rect 378 12928 3598 12968
rect 250 12068 314 12074
rect 380 12924 3598 12928
rect 380 12660 438 12924
rect 540 12890 606 12896
rect 540 12692 546 12890
rect 600 12692 606 12890
rect 540 12688 606 12692
rect 708 12660 754 12924
rect 856 12890 922 12896
rect 856 12692 862 12890
rect 916 12692 922 12890
rect 856 12688 922 12692
rect 1024 12660 1070 12924
rect 1172 12890 1238 12896
rect 1172 12692 1178 12890
rect 1232 12692 1238 12890
rect 1172 12688 1238 12692
rect 1340 12660 1386 12924
rect 1488 12890 1554 12896
rect 1488 12692 1494 12890
rect 1548 12692 1554 12890
rect 1488 12688 1554 12692
rect 1656 12660 1702 12924
rect 1804 12890 1870 12896
rect 1804 12692 1810 12890
rect 1864 12692 1870 12890
rect 1804 12688 1870 12692
rect 1972 12660 2018 12924
rect 2120 12890 2186 12896
rect 2120 12692 2126 12890
rect 2180 12692 2186 12890
rect 2120 12688 2186 12692
rect 2288 12660 2334 12924
rect 2436 12890 2502 12896
rect 2436 12692 2442 12890
rect 2496 12692 2502 12890
rect 2436 12688 2502 12692
rect 2604 12660 2650 12924
rect 2752 12890 2818 12896
rect 2752 12692 2758 12890
rect 2812 12692 2818 12890
rect 2752 12688 2818 12692
rect 2920 12660 2966 12924
rect 3068 12890 3134 12896
rect 3068 12692 3074 12890
rect 3128 12692 3134 12890
rect 3068 12688 3134 12692
rect 3236 12660 3282 12924
rect 3384 12890 3450 12896
rect 3384 12692 3390 12890
rect 3444 12692 3450 12890
rect 3384 12688 3450 12692
rect 3550 12660 3598 12924
rect 380 12614 3598 12660
rect 380 12350 438 12614
rect 540 12578 606 12582
rect 540 12386 546 12578
rect 600 12386 606 12578
rect 540 12382 606 12386
rect 708 12350 754 12614
rect 856 12578 922 12582
rect 856 12386 862 12578
rect 916 12386 922 12578
rect 856 12382 922 12386
rect 1024 12350 1070 12614
rect 1172 12578 1238 12582
rect 1172 12386 1178 12578
rect 1232 12386 1238 12578
rect 1172 12382 1238 12386
rect 1340 12350 1386 12614
rect 1488 12578 1554 12582
rect 1488 12386 1494 12578
rect 1548 12386 1554 12578
rect 1488 12382 1554 12386
rect 1656 12350 1702 12614
rect 1804 12578 1870 12582
rect 1804 12386 1810 12578
rect 1864 12386 1870 12578
rect 1804 12382 1870 12386
rect 1972 12350 2018 12614
rect 2120 12578 2186 12582
rect 2120 12386 2126 12578
rect 2180 12386 2186 12578
rect 2120 12382 2186 12386
rect 2288 12350 2334 12614
rect 2436 12578 2502 12582
rect 2436 12386 2442 12578
rect 2496 12386 2502 12578
rect 2436 12382 2502 12386
rect 2604 12350 2650 12614
rect 2752 12578 2818 12582
rect 2752 12386 2758 12578
rect 2812 12386 2818 12578
rect 2752 12382 2818 12386
rect 2920 12350 2966 12614
rect 3068 12578 3134 12582
rect 3068 12386 3074 12578
rect 3128 12386 3134 12578
rect 3068 12382 3134 12386
rect 3236 12350 3282 12614
rect 3384 12578 3450 12582
rect 3384 12386 3390 12578
rect 3444 12386 3450 12578
rect 3384 12382 3450 12386
rect 3550 12350 3598 12614
rect 380 12304 3598 12350
rect 380 12040 438 12304
rect 540 12268 606 12272
rect 540 12076 546 12268
rect 598 12076 606 12268
rect 540 12072 606 12076
rect 708 12040 754 12304
rect 856 12268 922 12272
rect 856 12076 862 12268
rect 914 12076 922 12268
rect 856 12072 922 12076
rect 1024 12040 1070 12304
rect 1172 12268 1238 12272
rect 1172 12076 1178 12268
rect 1230 12076 1238 12268
rect 1172 12072 1238 12076
rect 1340 12040 1386 12304
rect 1488 12268 1554 12272
rect 1488 12076 1494 12268
rect 1546 12076 1554 12268
rect 1488 12072 1554 12076
rect 1656 12040 1702 12304
rect 1804 12268 1870 12272
rect 1804 12076 1810 12268
rect 1862 12076 1870 12268
rect 1804 12072 1870 12076
rect 1972 12040 2018 12304
rect 2120 12268 2186 12272
rect 2120 12076 2126 12268
rect 2178 12076 2186 12268
rect 2120 12072 2186 12076
rect 2288 12040 2334 12304
rect 2436 12268 2502 12272
rect 2436 12076 2442 12268
rect 2494 12076 2502 12268
rect 2436 12072 2502 12076
rect 2604 12040 2650 12304
rect 2752 12268 2818 12272
rect 2752 12076 2758 12268
rect 2810 12076 2818 12268
rect 2752 12072 2818 12076
rect 2920 12040 2966 12304
rect 3068 12268 3134 12272
rect 3068 12076 3074 12268
rect 3126 12076 3134 12268
rect 3068 12072 3134 12076
rect 3236 12040 3282 12304
rect 3384 12268 3450 12272
rect 3384 12076 3390 12268
rect 3442 12076 3450 12268
rect 3384 12072 3450 12076
rect 3550 12040 3598 12304
rect 3676 12074 3692 13316
rect 3726 12074 3740 13316
rect 3676 12068 3740 12074
rect 380 11994 3598 12040
rect 380 11962 438 11994
rect 34 11730 438 11962
rect 540 11958 606 11962
rect 540 11766 546 11958
rect 598 11766 606 11958
rect 540 11762 606 11766
rect 708 11730 754 11994
rect 856 11958 922 11962
rect 856 11766 862 11958
rect 914 11766 922 11958
rect 856 11762 922 11766
rect 1024 11730 1070 11994
rect 1172 11958 1238 11962
rect 1172 11766 1178 11958
rect 1230 11766 1238 11958
rect 1172 11762 1238 11766
rect 1340 11730 1386 11994
rect 1488 11958 1554 11962
rect 1488 11766 1494 11958
rect 1546 11766 1554 11958
rect 1488 11762 1554 11766
rect 1656 11730 1702 11994
rect 1804 11958 1870 11962
rect 1804 11766 1810 11958
rect 1862 11766 1870 11958
rect 1804 11762 1870 11766
rect 1972 11730 2018 11994
rect 2120 11958 2186 11962
rect 2120 11766 2126 11958
rect 2178 11766 2186 11958
rect 2120 11762 2186 11766
rect 2288 11730 2334 11994
rect 2436 11958 2502 11962
rect 2436 11766 2442 11958
rect 2494 11766 2502 11958
rect 2436 11762 2502 11766
rect 2604 11730 2650 11994
rect 2752 11958 2818 11962
rect 2752 11766 2758 11958
rect 2810 11766 2818 11958
rect 2752 11762 2818 11766
rect 2920 11730 2966 11994
rect 3068 11958 3134 11962
rect 3068 11766 3074 11958
rect 3126 11766 3134 11958
rect 3068 11762 3134 11766
rect 3236 11730 3282 11994
rect 3550 11962 3598 11994
rect 3798 11962 4398 22106
rect 69346 13822 69954 13906
rect 69346 13324 69410 13822
rect 69866 13686 69954 13822
rect 70626 13686 70826 25646
rect 69866 13486 70826 13686
rect 69866 13324 69954 13486
rect 69346 13284 69954 13324
rect 3384 11958 3450 11962
rect 3384 11766 3390 11958
rect 3442 11766 3450 11958
rect 3384 11762 3450 11766
rect 3550 11730 4398 11962
rect -7122 11676 -3060 11694
rect -11792 11568 -11580 11574
rect -12162 11332 -11960 11348
rect -12162 10956 -12146 11332
rect -11974 11317 -11960 11332
rect -11974 10971 -11959 11317
rect -11974 10956 -11960 10971
rect -12162 10942 -11960 10956
rect -11792 10854 -11786 11568
rect -11586 10854 -11580 11568
rect -10386 11568 -10174 11574
rect -10756 11332 -10554 11348
rect -10756 10956 -10740 11332
rect -10568 11317 -10554 11332
rect -10568 10971 -10553 11317
rect -10568 10956 -10554 10971
rect -10756 10942 -10554 10956
rect -11792 10714 -11580 10854
rect -10386 10854 -10380 11568
rect -10180 10854 -10174 11568
rect -8980 11568 -8768 11574
rect -9350 11332 -9148 11348
rect -9350 10956 -9334 11332
rect -9162 11317 -9148 11332
rect -9162 10971 -9147 11317
rect -9162 10956 -9148 10971
rect -9350 10942 -9148 10956
rect -10386 10714 -10174 10854
rect -8980 10854 -8974 11568
rect -8774 10854 -8768 11568
rect -7574 11568 -7362 11574
rect -7944 11332 -7742 11348
rect -7944 10956 -7928 11332
rect -7756 11317 -7742 11332
rect -7756 10971 -7741 11317
rect -7756 10956 -7742 10971
rect -7944 10942 -7742 10956
rect -8980 10714 -8768 10854
rect -7574 10854 -7568 11568
rect -7368 10854 -7362 11568
rect -7122 11494 -3880 11676
rect -7574 10714 -7362 10854
rect -6744 11094 -3880 11494
rect -3280 11094 -3060 11676
rect 34 11684 4398 11730
rect 34 11452 438 11684
rect 540 11644 606 11652
rect 540 11456 546 11644
rect 598 11456 606 11644
rect 540 11452 606 11456
rect 380 11420 438 11452
rect 708 11420 754 11684
rect 856 11644 922 11652
rect 856 11456 862 11644
rect 914 11456 922 11644
rect 856 11452 922 11456
rect 1024 11420 1070 11684
rect 1172 11644 1238 11652
rect 1172 11456 1178 11644
rect 1230 11456 1238 11644
rect 1172 11452 1238 11456
rect 1340 11420 1386 11684
rect 1488 11644 1554 11652
rect 1488 11456 1494 11644
rect 1546 11456 1554 11644
rect 1488 11452 1554 11456
rect 1656 11420 1702 11684
rect 1804 11644 1870 11652
rect 1804 11456 1810 11644
rect 1862 11456 1870 11644
rect 1804 11452 1870 11456
rect 1972 11420 2018 11684
rect 2120 11644 2186 11652
rect 2120 11456 2126 11644
rect 2178 11456 2186 11644
rect 2120 11452 2186 11456
rect 2288 11420 2334 11684
rect 2436 11644 2502 11652
rect 2436 11456 2442 11644
rect 2494 11456 2502 11644
rect 2436 11452 2502 11456
rect 2604 11420 2650 11684
rect 2752 11644 2818 11652
rect 2752 11456 2758 11644
rect 2810 11456 2818 11644
rect 2752 11452 2818 11456
rect 2920 11420 2966 11684
rect 3068 11644 3134 11652
rect 3068 11456 3074 11644
rect 3126 11456 3134 11644
rect 3068 11452 3134 11456
rect 3236 11420 3282 11684
rect 3384 11644 3450 11652
rect 3384 11456 3390 11644
rect 3442 11456 3450 11644
rect 3384 11452 3450 11456
rect 3550 11452 4398 11684
rect 3550 11420 3598 11452
rect 380 11374 3598 11420
rect 250 11340 314 11346
rect -6744 10694 -6144 11094
rect -7122 10494 -6144 10694
rect -11792 9962 -11580 9968
rect -12162 9726 -11960 9742
rect -12162 9350 -12146 9726
rect -11974 9711 -11960 9726
rect -11974 9365 -11959 9711
rect -11974 9350 -11960 9365
rect -12162 9336 -11960 9350
rect -11792 9114 -11786 9962
rect -11586 9114 -11580 9962
rect -10386 9962 -10174 9968
rect -10756 9726 -10554 9742
rect -10756 9350 -10740 9726
rect -10568 9711 -10554 9726
rect -10568 9365 -10553 9711
rect -10568 9350 -10554 9365
rect -10756 9336 -10554 9350
rect -11792 9108 -11580 9114
rect -10386 9114 -10380 9962
rect -10180 9114 -10174 9962
rect -8980 9962 -8768 9968
rect -9350 9726 -9148 9742
rect -9350 9350 -9334 9726
rect -9162 9711 -9148 9726
rect -9162 9365 -9147 9711
rect -9162 9350 -9148 9365
rect -9350 9336 -9148 9350
rect -10386 9108 -10174 9114
rect -8980 9114 -8974 9962
rect -8774 9114 -8768 9962
rect -7574 9962 -7362 9968
rect -7944 9726 -7742 9742
rect -7944 9350 -7928 9726
rect -7756 9711 -7742 9726
rect -7756 9365 -7741 9711
rect -7756 9350 -7742 9365
rect -7944 9336 -7742 9350
rect -8980 9108 -8768 9114
rect -7574 9114 -7568 9962
rect -7368 9114 -7362 9962
rect -6744 9906 -6144 10494
rect 250 10098 264 11340
rect 298 10098 314 11340
rect 380 11110 438 11374
rect 540 11334 606 11342
rect 540 11146 546 11334
rect 598 11146 606 11334
rect 540 11142 606 11146
rect 708 11110 754 11374
rect 856 11334 922 11342
rect 856 11146 862 11334
rect 914 11146 922 11334
rect 856 11142 922 11146
rect 1024 11110 1070 11374
rect 1172 11334 1238 11342
rect 1172 11146 1178 11334
rect 1230 11146 1238 11334
rect 1172 11142 1238 11146
rect 1340 11110 1386 11374
rect 1488 11334 1554 11342
rect 1488 11146 1494 11334
rect 1546 11146 1554 11334
rect 1488 11142 1554 11146
rect 1656 11110 1702 11374
rect 1804 11334 1870 11342
rect 1804 11146 1810 11334
rect 1862 11146 1870 11334
rect 1804 11142 1870 11146
rect 1972 11110 2018 11374
rect 2120 11334 2186 11342
rect 2120 11146 2126 11334
rect 2178 11146 2186 11334
rect 2120 11142 2186 11146
rect 2288 11110 2334 11374
rect 2436 11334 2502 11342
rect 2436 11146 2442 11334
rect 2494 11146 2502 11334
rect 2436 11142 2502 11146
rect 2604 11110 2650 11374
rect 2752 11334 2818 11342
rect 2752 11146 2758 11334
rect 2810 11146 2818 11334
rect 2752 11142 2818 11146
rect 2920 11110 2966 11374
rect 3068 11334 3134 11342
rect 3068 11146 3074 11334
rect 3126 11146 3134 11334
rect 3068 11142 3134 11146
rect 3236 11110 3282 11374
rect 3384 11334 3450 11342
rect 3384 11146 3390 11334
rect 3442 11146 3450 11334
rect 3384 11142 3450 11146
rect 3550 11110 3598 11374
rect 380 11064 3598 11110
rect 380 10800 438 11064
rect 540 11026 606 11032
rect 540 10838 546 11026
rect 598 10838 606 11026
rect 540 10832 606 10838
rect 708 10800 754 11064
rect 856 11026 922 11032
rect 856 10838 862 11026
rect 914 10838 922 11026
rect 856 10832 922 10838
rect 1024 10800 1070 11064
rect 1172 11026 1238 11032
rect 1172 10838 1178 11026
rect 1230 10838 1238 11026
rect 1172 10832 1238 10838
rect 1340 10800 1386 11064
rect 1488 11026 1554 11032
rect 1488 10838 1494 11026
rect 1546 10838 1554 11026
rect 1488 10832 1554 10838
rect 1656 10800 1702 11064
rect 1804 11026 1870 11032
rect 1804 10838 1810 11026
rect 1862 10838 1870 11026
rect 1804 10832 1870 10838
rect 1972 10800 2018 11064
rect 2120 11026 2186 11032
rect 2120 10838 2126 11026
rect 2178 10838 2186 11026
rect 2120 10832 2186 10838
rect 2288 10800 2334 11064
rect 2436 11026 2502 11032
rect 2436 10838 2442 11026
rect 2494 10838 2502 11026
rect 2436 10832 2502 10838
rect 2604 10800 2650 11064
rect 2752 11026 2818 11032
rect 2752 10838 2758 11026
rect 2810 10838 2818 11026
rect 2752 10832 2818 10838
rect 2920 10800 2966 11064
rect 3068 11026 3134 11032
rect 3068 10838 3074 11026
rect 3126 10838 3134 11026
rect 3068 10832 3134 10838
rect 3236 10800 3282 11064
rect 3384 11026 3450 11032
rect 3384 10838 3390 11026
rect 3442 10838 3450 11026
rect 3384 10832 3450 10838
rect 3550 10800 3598 11064
rect 380 10754 3598 10800
rect 380 10490 438 10754
rect 540 10712 606 10722
rect 540 10526 546 10712
rect 598 10526 606 10712
rect 540 10522 606 10526
rect 708 10490 754 10754
rect 856 10712 922 10722
rect 856 10526 862 10712
rect 914 10526 922 10712
rect 856 10522 922 10526
rect 1024 10490 1070 10754
rect 1172 10712 1238 10722
rect 1172 10526 1178 10712
rect 1230 10526 1238 10712
rect 1172 10522 1238 10526
rect 1340 10490 1386 10754
rect 1488 10712 1554 10722
rect 1488 10526 1494 10712
rect 1546 10526 1554 10712
rect 1488 10522 1554 10526
rect 1656 10490 1702 10754
rect 1804 10712 1870 10722
rect 1804 10526 1810 10712
rect 1862 10526 1870 10712
rect 1804 10522 1870 10526
rect 1972 10490 2018 10754
rect 2120 10712 2186 10722
rect 2120 10526 2126 10712
rect 2178 10526 2186 10712
rect 2120 10522 2186 10526
rect 2288 10490 2334 10754
rect 2436 10712 2502 10722
rect 2436 10526 2442 10712
rect 2494 10526 2502 10712
rect 2436 10522 2502 10526
rect 2604 10490 2650 10754
rect 2752 10712 2818 10722
rect 2752 10526 2758 10712
rect 2810 10526 2818 10712
rect 2752 10522 2818 10526
rect 2920 10490 2966 10754
rect 3068 10712 3134 10722
rect 3068 10526 3074 10712
rect 3126 10526 3134 10712
rect 3068 10522 3134 10526
rect 3236 10490 3282 10754
rect 3384 10712 3450 10722
rect 3384 10526 3390 10712
rect 3442 10526 3450 10712
rect 3384 10522 3450 10526
rect 3550 10490 3598 10754
rect 380 10444 3598 10490
rect 380 10180 438 10444
rect 540 10404 606 10412
rect 540 10218 546 10404
rect 598 10218 606 10404
rect 540 10208 606 10218
rect 708 10180 754 10444
rect 856 10404 922 10412
rect 856 10218 862 10404
rect 914 10218 922 10404
rect 856 10208 922 10218
rect 1024 10180 1070 10444
rect 1172 10404 1238 10412
rect 1172 10218 1178 10404
rect 1230 10218 1238 10404
rect 1172 10208 1238 10218
rect 1340 10180 1386 10444
rect 1488 10404 1554 10412
rect 1488 10218 1494 10404
rect 1546 10218 1554 10404
rect 1488 10208 1554 10218
rect 1656 10180 1702 10444
rect 1804 10404 1870 10412
rect 1804 10218 1810 10404
rect 1862 10218 1870 10404
rect 1804 10208 1870 10218
rect 1972 10180 2018 10444
rect 2120 10404 2186 10412
rect 2120 10218 2126 10404
rect 2178 10218 2186 10404
rect 2120 10208 2186 10218
rect 2288 10180 2334 10444
rect 2436 10404 2502 10412
rect 2436 10218 2442 10404
rect 2494 10218 2502 10404
rect 2436 10208 2502 10218
rect 2604 10180 2650 10444
rect 2752 10404 2818 10412
rect 2752 10218 2758 10404
rect 2810 10218 2818 10404
rect 2752 10208 2818 10218
rect 2920 10180 2966 10444
rect 3068 10404 3134 10412
rect 3068 10218 3074 10404
rect 3126 10218 3134 10404
rect 3068 10208 3134 10218
rect 3236 10180 3282 10444
rect 3384 10404 3450 10412
rect 3384 10218 3390 10404
rect 3442 10218 3450 10404
rect 3384 10208 3450 10218
rect 3550 10180 3598 10444
rect 380 10120 3598 10180
rect 3678 11340 3742 11346
rect 250 10052 314 10098
rect 3678 10098 3692 11340
rect 3726 10098 3742 11340
rect 3678 10052 3742 10098
rect 250 10046 3742 10052
rect 250 10036 544 10046
rect 250 10002 360 10036
rect 3446 10036 3742 10046
rect 3630 10002 3742 10036
rect 250 9994 544 10002
rect 3446 9994 3742 10002
rect 250 9988 3742 9994
rect -6744 9706 -4760 9906
rect -6744 9694 -6144 9706
rect -7122 9494 -6144 9694
rect -4164 9494 -3964 9894
rect -7574 9108 -7362 9114
rect -6744 8694 -6144 9494
rect -4778 8988 -4378 9188
rect -3768 8984 -3368 9184
rect -7122 8494 -6144 8694
rect -6744 8442 -6144 8494
rect -11792 8356 -11580 8362
rect -12162 8120 -11960 8136
rect -12162 7744 -12146 8120
rect -11974 7744 -11960 8120
rect -12162 7730 -11960 7744
rect -11792 7508 -11786 8356
rect -11586 7508 -11580 8356
rect -10386 8356 -10174 8362
rect -10756 8120 -10554 8136
rect -10756 7744 -10740 8120
rect -10568 8105 -10554 8120
rect -10568 7759 -10553 8105
rect -10568 7744 -10554 7759
rect -10756 7730 -10554 7744
rect -11792 7502 -11580 7508
rect -10386 7508 -10380 8356
rect -10180 7508 -10174 8356
rect -8980 8356 -8768 8362
rect -9350 8120 -9148 8136
rect -9350 7744 -9334 8120
rect -9162 8105 -9148 8120
rect -9162 7759 -9147 8105
rect -9162 7744 -9148 7759
rect -9350 7730 -9148 7744
rect -10386 7502 -10174 7508
rect -8980 7508 -8974 8356
rect -8774 7508 -8768 8356
rect -7574 8356 -7362 8362
rect -7944 8120 -7742 8136
rect -7944 7744 -7928 8120
rect -7756 8105 -7742 8120
rect -7756 7759 -7741 8105
rect -7756 7744 -7742 7759
rect -7944 7730 -7742 7744
rect -8980 7502 -8768 7508
rect -7574 7508 -7568 8356
rect -7368 7508 -7362 8356
rect -6744 8242 -4776 8442
rect -4160 8262 -3960 8662
rect -6744 7694 -6144 8242
rect -7574 7502 -7362 7508
rect -7122 7494 -6144 7694
rect -11792 6750 -11580 6756
rect -12162 6514 -11960 6530
rect -12162 6138 -12146 6514
rect -11974 6138 -11960 6514
rect -12162 6124 -11960 6138
rect -11792 5902 -11786 6750
rect -11586 5902 -11580 6750
rect -10386 6750 -10174 6756
rect -10756 6514 -10554 6530
rect -10756 6138 -10740 6514
rect -10568 6499 -10554 6514
rect -10568 6153 -10553 6499
rect -10568 6138 -10554 6153
rect -10756 6124 -10554 6138
rect -11792 5896 -11580 5902
rect -10386 5902 -10380 6750
rect -10180 5902 -10174 6750
rect -8980 6750 -8768 6756
rect -9350 6514 -9148 6530
rect -9350 6138 -9334 6514
rect -9162 6499 -9148 6514
rect -9162 6153 -9147 6499
rect -9162 6138 -9148 6153
rect -9350 6124 -9148 6138
rect -10386 5896 -10174 5902
rect -8980 5902 -8974 6750
rect -8774 5902 -8768 6750
rect -7574 6750 -7362 6756
rect -7944 6514 -7742 6530
rect -7944 6138 -7928 6514
rect -7756 6499 -7742 6514
rect -7756 6153 -7741 6499
rect -7756 6138 -7742 6153
rect -7944 6124 -7742 6138
rect -8980 5896 -8768 5902
rect -7574 5902 -7568 6750
rect -7368 5902 -7362 6750
rect -6744 6694 -6144 7494
rect -7122 6494 -6144 6694
rect -7574 5896 -7362 5902
rect -6744 5998 -6144 6494
rect -6744 5694 -6148 5998
rect -7122 5494 -6148 5694
<< via1 >>
rect -1522 30310 7242 30854
rect -1522 30276 -1358 30310
rect -1358 30276 -310 30310
rect -310 30276 38 30310
rect 38 30276 1086 30310
rect 1086 30276 1434 30310
rect 1434 30276 2482 30310
rect 2482 30276 2830 30310
rect 2830 30276 3878 30310
rect 3878 30276 7242 30310
rect -1522 30274 7242 30276
rect -17786 28472 -17590 28872
rect -17404 28254 -17222 29096
rect -16380 28472 -16184 28872
rect -15998 28254 -15816 29096
rect -14974 28472 -14778 28872
rect -14592 28254 -14410 29096
rect -13568 28472 -13372 28872
rect -13186 28254 -13004 29096
rect -12162 28472 -11966 28872
rect -11780 28254 -11598 29096
rect -10756 28472 -10560 28872
rect -10374 28254 -10192 29096
rect -9350 28472 -9154 28872
rect -8968 28254 -8786 29096
rect -7944 28472 -7748 28872
rect -7562 28254 -7380 29096
rect -6538 28472 -6342 28872
rect -6156 28254 -5974 29096
rect -5132 28472 -4936 28872
rect -4750 28254 -4568 29096
rect -17786 26866 -17590 27266
rect -17404 26648 -17222 27490
rect -16380 26866 -16184 27266
rect -15998 26648 -15816 27490
rect -14974 26866 -14778 27266
rect -14592 26648 -14410 27490
rect -13568 26866 -13372 27266
rect -13186 26648 -13004 27490
rect -12162 26866 -11966 27266
rect -11780 26648 -11598 27490
rect -10756 26866 -10560 27266
rect -10374 26648 -10192 27490
rect -9350 26866 -9154 27266
rect -8968 26648 -8786 27490
rect -7944 26866 -7748 27266
rect -7562 26648 -7380 27490
rect -6538 26866 -6342 27266
rect -6156 26648 -5974 27490
rect -5132 26866 -4936 27266
rect -4750 26648 -4568 27490
rect -17786 25260 -17590 25660
rect -17404 25042 -17222 25884
rect -16380 25260 -16184 25660
rect -15998 25042 -15816 25884
rect -14974 25260 -14778 25660
rect -14592 25042 -14410 25884
rect -13568 25260 -13372 25660
rect -13186 25042 -13004 25884
rect -12162 25260 -11966 25660
rect -11780 25042 -11598 25884
rect -10756 25260 -10560 25660
rect -10374 25042 -10192 25884
rect -9350 25260 -9154 25660
rect -8968 25042 -8786 25884
rect -7944 25260 -7748 25660
rect -7562 25042 -7380 25884
rect -6538 25260 -6342 25660
rect -6156 25042 -5974 25884
rect -5132 25260 -4936 25660
rect -4750 25042 -4568 25884
rect -2982 24656 -2396 30034
rect -1224 29300 -444 30080
rect 172 29300 952 30080
rect 1568 29300 2348 30080
rect 2964 29300 3744 30080
rect -1696 28878 -1368 29106
rect -300 28878 28 29106
rect 1096 28878 1424 29106
rect 2492 28878 2820 29106
rect 3888 28878 4216 29106
rect -1224 27904 -444 28684
rect 172 27904 952 28684
rect 1568 27904 2348 28684
rect 2964 27904 3744 28684
rect -1696 27482 -1368 27710
rect -300 27482 28 27710
rect 1096 27482 1424 27710
rect 2492 27482 2820 27710
rect 3888 27482 4216 27710
rect -1224 26508 -444 27288
rect 172 26508 952 27288
rect 1568 26508 2348 27288
rect 2964 26508 3744 27288
rect -1696 26086 -1368 26314
rect -300 26086 28 26314
rect 1096 26086 1424 26314
rect 2492 26086 2820 26314
rect 3888 26086 4216 26314
rect -1224 25112 -444 25892
rect 172 25112 952 25892
rect 1568 25112 2348 25892
rect 2964 25112 3744 25892
rect 9820 27342 10600 28122
rect 10796 27208 10830 28256
rect 10830 27208 10986 28256
rect 10986 27208 11020 28256
rect 9820 25946 10600 26726
rect 10796 26860 11020 27208
rect 11216 27342 11996 28122
rect 12192 27208 12226 28256
rect 12226 27208 12382 28256
rect 12382 27208 12416 28256
rect 10796 25812 10830 26860
rect 10830 25812 10986 26860
rect 10986 25812 11020 26860
rect 10796 25716 11020 25812
rect 11216 25946 11996 26726
rect 12192 26860 12416 27208
rect 12612 27342 13392 28122
rect 13588 27208 13622 28256
rect 13622 27208 13778 28256
rect 13778 27208 13812 28256
rect 12192 25812 12226 26860
rect 12226 25812 12382 26860
rect 12382 25812 12416 26860
rect 12192 25716 12416 25812
rect 12612 25946 13392 26726
rect 13588 26860 13812 27208
rect 14008 27342 14788 28122
rect 14984 27208 15018 28256
rect 15018 27208 15174 28256
rect 15174 27208 15208 28256
rect 13588 25812 13622 26860
rect 13622 25812 13778 26860
rect 13778 25812 13812 26860
rect 13588 25716 13812 25812
rect 14008 25946 14788 26726
rect 14984 26860 15208 27208
rect 15404 27342 16184 28122
rect 16380 27208 16414 28256
rect 16414 27208 16570 28256
rect 16570 27208 16604 28256
rect 14984 25812 15018 26860
rect 15018 25812 15174 26860
rect 15174 25812 15208 26860
rect 14984 25716 15208 25812
rect 15404 25946 16184 26726
rect 16380 26860 16604 27208
rect 16800 27342 17580 28122
rect 17776 27208 17810 28256
rect 17810 27208 17966 28256
rect 17966 27208 18000 28256
rect 16380 25812 16414 26860
rect 16414 25812 16570 26860
rect 16570 25812 16604 26860
rect 16380 25716 16604 25812
rect 16800 25946 17580 26726
rect 17776 26860 18000 27208
rect 18196 27342 18976 28122
rect 19172 27208 19206 28256
rect 19206 27208 19362 28256
rect 19362 27208 19396 28256
rect 17776 25812 17810 26860
rect 17810 25812 17966 26860
rect 17966 25812 18000 26860
rect 17776 25716 18000 25812
rect 18196 25946 18976 26726
rect 19172 26860 19396 27208
rect 19592 27342 20372 28122
rect 20568 27208 20602 28256
rect 20602 27208 20758 28256
rect 20758 27208 20792 28256
rect 19172 25812 19206 26860
rect 19206 25812 19362 26860
rect 19362 25812 19396 26860
rect 19172 25716 19396 25812
rect 19592 25946 20372 26726
rect 20568 26860 20792 27208
rect 20988 27342 21768 28122
rect 21964 27208 21998 28256
rect 21998 27208 22154 28256
rect 22154 27208 22188 28256
rect 20568 25812 20602 26860
rect 20602 25812 20758 26860
rect 20758 25812 20792 26860
rect 20568 25716 20792 25812
rect 20988 25946 21768 26726
rect 21964 26860 22188 27208
rect 22384 27342 23164 28122
rect 23360 27208 23394 28256
rect 23394 27208 23550 28256
rect 23550 27208 23584 28256
rect 21964 25812 21998 26860
rect 21998 25812 22154 26860
rect 22154 25812 22188 26860
rect 21964 25716 22188 25812
rect 22384 25946 23164 26726
rect 23360 26860 23584 27208
rect 23780 27342 24560 28122
rect 24756 27208 24790 28256
rect 24790 27208 24946 28256
rect 24946 27208 24980 28256
rect 23360 25812 23394 26860
rect 23394 25812 23550 26860
rect 23550 25812 23584 26860
rect 23360 25716 23584 25812
rect 23780 25946 24560 26726
rect 24756 26860 24980 27208
rect 25176 27342 25956 28122
rect 26152 27208 26186 28256
rect 26186 27208 26342 28256
rect 26342 27208 26376 28256
rect 24756 25812 24790 26860
rect 24790 25812 24946 26860
rect 24946 25812 24980 26860
rect 24756 25716 24980 25812
rect 25176 25946 25956 26726
rect 26152 26860 26376 27208
rect 26572 27342 27352 28122
rect 27548 27208 27582 28256
rect 27582 27208 27738 28256
rect 27738 27208 27772 28256
rect 26152 25812 26186 26860
rect 26186 25812 26342 26860
rect 26342 25812 26376 26860
rect 26152 25716 26376 25812
rect 26572 25946 27352 26726
rect 27548 26860 27772 27208
rect 27968 27342 28748 28122
rect 28944 27208 28978 28256
rect 28978 27208 29134 28256
rect 29134 27208 29168 28256
rect 27548 25812 27582 26860
rect 27582 25812 27738 26860
rect 27738 25812 27772 26860
rect 27548 25716 27772 25812
rect 27968 25946 28748 26726
rect 28944 26860 29168 27208
rect 29362 27342 30144 28122
rect 30340 27208 30374 28256
rect 30374 27208 30530 28256
rect 30530 27208 30564 28256
rect 28944 25812 28978 26860
rect 28978 25812 29134 26860
rect 29134 25812 29168 26860
rect 28944 25716 29168 25812
rect 29362 25946 30144 26726
rect 30340 26860 30564 27208
rect 30760 27342 31540 28122
rect 31736 27208 31770 28256
rect 31770 27208 31926 28256
rect 31926 27208 31960 28256
rect 30340 25812 30374 26860
rect 30374 25812 30530 26860
rect 30530 25812 30564 26860
rect 30340 25716 30564 25812
rect 30760 25946 31540 26726
rect 31736 26860 31960 27208
rect 32156 27342 32936 28122
rect 33132 27208 33166 28256
rect 33166 27208 33322 28256
rect 33322 27208 33356 28256
rect 31736 25812 31770 26860
rect 31770 25812 31926 26860
rect 31926 25812 31960 26860
rect 31736 25716 31960 25812
rect 32156 25946 32936 26726
rect 33132 26860 33356 27208
rect 33552 27342 34332 28122
rect 34528 27208 34562 28256
rect 34562 27208 34718 28256
rect 34718 27208 34752 28256
rect 33132 25812 33166 26860
rect 33166 25812 33322 26860
rect 33322 25812 33356 26860
rect 33132 25716 33356 25812
rect 33552 25946 34332 26726
rect 34528 26860 34752 27208
rect 34948 27342 35728 28122
rect 35924 27208 35958 28256
rect 35958 27208 36114 28256
rect 36114 27208 36148 28256
rect 34528 25812 34562 26860
rect 34562 25812 34718 26860
rect 34718 25812 34752 26860
rect 34528 25716 34752 25812
rect 34948 25946 35728 26726
rect 35924 26860 36148 27208
rect 36344 27342 37124 28122
rect 37320 27208 37354 28256
rect 37354 27208 37510 28256
rect 37510 27208 37544 28256
rect 35924 25812 35958 26860
rect 35958 25812 36114 26860
rect 36114 25812 36148 26860
rect 35924 25716 36148 25812
rect 36344 25946 37124 26726
rect 37320 26860 37544 27208
rect 37740 27342 38520 28122
rect 38716 27208 38750 28256
rect 38750 27208 38906 28256
rect 38906 27208 38940 28256
rect 37320 25812 37354 26860
rect 37354 25812 37510 26860
rect 37510 25812 37544 26860
rect 37320 25716 37544 25812
rect 37740 25946 38520 26726
rect 38716 26860 38940 27208
rect 39136 27342 39916 28122
rect 40112 27208 40146 28256
rect 40146 27208 40302 28256
rect 40302 27208 40336 28256
rect 38716 25812 38750 26860
rect 38750 25812 38906 26860
rect 38906 25812 38940 26860
rect 38716 25716 38940 25812
rect 39136 25946 39916 26726
rect 40112 26860 40336 27208
rect 40532 27342 41312 28122
rect 41508 27208 41542 28256
rect 41542 27208 41698 28256
rect 41698 27208 41732 28256
rect 40112 25812 40146 26860
rect 40146 25812 40302 26860
rect 40302 25812 40336 26860
rect 40112 25716 40336 25812
rect 40532 25946 41312 26726
rect 41508 26860 41732 27208
rect 41928 27342 42708 28122
rect 42904 27208 42938 28256
rect 42938 27208 43094 28256
rect 43094 27208 43128 28256
rect 41508 25812 41542 26860
rect 41542 25812 41698 26860
rect 41698 25812 41732 26860
rect 41508 25716 41732 25812
rect 41928 25946 42708 26726
rect 42904 26860 43128 27208
rect 43324 27342 44104 28122
rect 44300 27208 44334 28256
rect 44334 27208 44490 28256
rect 44490 27208 44524 28256
rect 42904 25812 42938 26860
rect 42938 25812 43094 26860
rect 43094 25812 43128 26860
rect 42904 25716 43128 25812
rect 43324 25946 44104 26726
rect 44300 26860 44524 27208
rect 44720 27342 45500 28122
rect 45696 27208 45730 28256
rect 45730 27208 45886 28256
rect 45886 27208 45920 28256
rect 44300 25812 44334 26860
rect 44334 25812 44490 26860
rect 44490 25812 44524 26860
rect 44300 25716 44524 25812
rect 44720 25946 45500 26726
rect 45696 26860 45920 27208
rect 46116 27342 46896 28122
rect 47092 27208 47126 28256
rect 47126 27208 47282 28256
rect 47282 27208 47316 28256
rect 45696 25812 45730 26860
rect 45730 25812 45886 26860
rect 45886 25812 45920 26860
rect 45696 25716 45920 25812
rect 46116 25946 46896 26726
rect 47092 26860 47316 27208
rect 47512 27342 48292 28122
rect 48488 27208 48522 28256
rect 48522 27208 48678 28256
rect 48678 27208 48712 28256
rect 47092 25812 47126 26860
rect 47126 25812 47282 26860
rect 47282 25812 47316 26860
rect 47092 25716 47316 25812
rect 47512 25946 48292 26726
rect 48488 26860 48712 27208
rect 48908 27342 49688 28122
rect 49884 27208 49918 28256
rect 49918 27208 50074 28256
rect 50074 27208 50108 28256
rect 48488 25812 48522 26860
rect 48522 25812 48678 26860
rect 48678 25812 48712 26860
rect 48488 25716 48712 25812
rect 48908 25946 49688 26726
rect 49884 26860 50108 27208
rect 50304 27342 51084 28122
rect 49884 25812 49918 26860
rect 49918 25812 50074 26860
rect 50074 25812 50108 26860
rect 49884 25716 50108 25812
rect 50304 25946 51084 26726
rect -1696 24690 -1368 24918
rect -300 24690 28 24918
rect 1096 24690 1424 24918
rect 2492 24690 2820 24918
rect 3888 24690 4216 24918
rect -17786 23654 -17590 24054
rect -17404 23436 -17222 24278
rect -16380 23654 -16184 24054
rect -15998 23436 -15816 24278
rect -14974 23654 -14778 24054
rect -14592 23436 -14410 24278
rect -13568 23654 -13372 24054
rect -13186 23436 -13004 24278
rect -12162 23654 -11966 24054
rect -11780 23436 -11598 24278
rect -10756 23654 -10560 24054
rect -10374 23436 -10192 24278
rect -9350 23654 -9154 24054
rect -8968 23436 -8786 24278
rect -7944 23654 -7748 24054
rect -7562 23436 -7380 24278
rect -6538 23654 -6342 24054
rect -6156 23436 -5974 24278
rect -5132 23654 -4936 24054
rect -4750 23436 -4568 24278
rect -1228 23856 3618 24438
rect -17786 22048 -17590 22448
rect -17404 21830 -17222 22672
rect -16380 22048 -16184 22448
rect -15998 21830 -15816 22672
rect -14974 22048 -14778 22448
rect -14592 21830 -14410 22672
rect -13568 22048 -13372 22448
rect -13186 21830 -13004 22672
rect -12162 22048 -11966 22448
rect -11780 21830 -11598 22672
rect -10756 22048 -10560 22448
rect -10374 21830 -10192 22672
rect -9350 22048 -9154 22448
rect -8968 21830 -8786 22672
rect -7944 22048 -7748 22448
rect -7562 21830 -7380 22672
rect -6538 22048 -6342 22448
rect -6156 21830 -5974 22672
rect -5132 22048 -4936 22448
rect -4750 21830 -4568 22672
rect -17786 20442 -17590 20842
rect -17404 20224 -17222 21066
rect -16380 20442 -16184 20842
rect -15998 20224 -15816 21066
rect -14974 20442 -14778 20842
rect -14592 20224 -14410 21066
rect -13568 20442 -13372 20842
rect -13186 20224 -13004 21066
rect -12162 20442 -11966 20842
rect -11780 20224 -11598 21066
rect -10756 20442 -10560 20842
rect -10374 20224 -10192 21066
rect -9350 20442 -9154 20842
rect -8968 20224 -8786 21066
rect -7944 20442 -7748 20842
rect -7562 20224 -7380 21066
rect -6538 20442 -6342 20842
rect -6156 20224 -5974 21066
rect -5132 20442 -4936 20842
rect -4750 20224 -4568 21066
rect 3698 22936 4098 23336
rect -17786 18836 -17590 19236
rect -17404 18618 -17222 19460
rect -16380 18836 -16184 19236
rect -15998 18618 -15816 19460
rect -14974 18836 -14778 19236
rect -14592 18618 -14410 19460
rect -13568 18836 -13372 19236
rect -13186 18618 -13004 19460
rect -12162 18836 -11966 19236
rect -11780 18618 -11598 19460
rect -10756 18836 -10560 19236
rect -10374 18618 -10192 19460
rect -9350 18836 -9154 19236
rect -8968 18618 -8786 19460
rect -7944 18836 -7748 19236
rect -7562 18618 -7380 19460
rect -6538 18836 -6342 19236
rect -6156 18618 -5974 19460
rect -5132 18836 -4936 19236
rect -4750 18618 -4568 19460
rect -2968 19016 -2568 19040
rect -2968 18664 -2944 19016
rect -2944 18664 -2592 19016
rect -2592 18664 -2568 19016
rect -2968 18640 -2568 18664
rect -17786 17230 -17590 17630
rect -17404 17012 -17222 17854
rect -16380 17230 -16184 17630
rect -15998 17012 -15816 17854
rect -14974 17230 -14778 17630
rect -14592 17012 -14410 17854
rect -13568 17230 -13372 17630
rect -13186 17012 -13004 17854
rect -12162 17230 -11966 17630
rect -11780 17012 -11598 17854
rect -10756 17230 -10560 17630
rect -10374 17012 -10192 17854
rect -9350 17230 -9154 17630
rect -8968 17012 -8786 17854
rect -7944 17230 -7748 17630
rect -7562 17012 -7380 17854
rect -6538 17230 -6342 17630
rect -6156 17012 -5974 17854
rect -5132 17230 -4936 17630
rect -4750 17012 -4568 17854
rect -17786 15624 -17590 16024
rect -17404 15406 -17222 16248
rect -16380 15624 -16184 16024
rect -15998 15406 -15816 16248
rect -14974 15624 -14778 16024
rect -14592 15406 -14410 16248
rect -13568 15624 -13372 16024
rect -13186 15406 -13004 16248
rect -12162 15624 -11966 16024
rect -11780 15406 -11598 16248
rect -10756 15624 -10560 16024
rect -10374 15406 -10192 16248
rect -9350 15624 -9154 16024
rect -8968 15406 -8786 16248
rect -7944 15624 -7748 16024
rect -7562 15406 -7380 16248
rect -6538 15624 -6342 16024
rect -6156 15406 -5974 16248
rect -5132 15624 -4936 16024
rect -4750 15406 -4568 16248
rect -17786 14018 -17590 14418
rect -17404 13800 -17222 14642
rect -16380 14018 -16184 14418
rect -15998 13800 -15816 14642
rect -14974 14018 -14778 14418
rect -14592 13800 -14410 14642
rect -13568 14018 -13372 14418
rect -13186 13800 -13004 14642
rect -12162 14018 -11966 14418
rect -11780 13800 -11598 14642
rect -10756 14018 -10560 14418
rect -10374 13800 -10192 14642
rect -9350 14018 -9154 14418
rect -8968 13800 -8786 14642
rect -7944 14018 -7748 14418
rect -7562 13800 -7380 14642
rect -6538 14018 -6342 14418
rect -6156 13800 -5974 14642
rect -5132 14018 -4936 14418
rect -4750 13800 -4568 14642
rect 538 13412 604 13426
rect 604 13412 3448 13426
rect 538 13378 3448 13412
rect 538 13370 604 13378
rect 604 13370 3448 13378
rect 546 13004 600 13202
rect 862 13004 916 13202
rect 1178 13004 1232 13202
rect 1494 13004 1548 13202
rect 1810 13004 1864 13202
rect 2126 13004 2180 13202
rect 2442 13004 2496 13202
rect 2758 13004 2812 13202
rect 3074 13004 3128 13202
rect 3390 13004 3444 13202
rect 546 12692 600 12890
rect 862 12692 916 12890
rect 1178 12692 1232 12890
rect 1494 12692 1548 12890
rect 1810 12692 1864 12890
rect 2126 12692 2180 12890
rect 2442 12692 2496 12890
rect 2758 12692 2812 12890
rect 3074 12692 3128 12890
rect 3390 12692 3444 12890
rect 546 12386 600 12578
rect 862 12386 916 12578
rect 1178 12386 1232 12578
rect 1494 12386 1548 12578
rect 1810 12386 1864 12578
rect 2126 12386 2180 12578
rect 2442 12386 2496 12578
rect 2758 12386 2812 12578
rect 3074 12386 3128 12578
rect 3390 12386 3444 12578
rect 546 12076 598 12268
rect 862 12076 914 12268
rect 1178 12076 1230 12268
rect 1494 12076 1546 12268
rect 1810 12076 1862 12268
rect 2126 12076 2178 12268
rect 2442 12076 2494 12268
rect 2758 12076 2810 12268
rect 3074 12076 3126 12268
rect 3390 12076 3442 12268
rect 546 11766 598 11958
rect 862 11766 914 11958
rect 1178 11766 1230 11958
rect 1494 11766 1546 11958
rect 1810 11766 1862 11958
rect 2126 11766 2178 11958
rect 2442 11766 2494 11958
rect 2758 11766 2810 11958
rect 3074 11766 3126 11958
rect 69410 13324 69866 13822
rect 3390 11766 3442 11958
rect -12146 10956 -11974 11332
rect -11786 10854 -11586 11568
rect -10740 10956 -10568 11332
rect -10380 10854 -10180 11568
rect -9334 10956 -9162 11332
rect -8974 10854 -8774 11568
rect -7928 10956 -7756 11332
rect -7568 10854 -7368 11568
rect -3880 11094 -3280 11676
rect 546 11456 598 11644
rect 862 11456 914 11644
rect 1178 11456 1230 11644
rect 1494 11456 1546 11644
rect 1810 11456 1862 11644
rect 2126 11456 2178 11644
rect 2442 11456 2494 11644
rect 2758 11456 2810 11644
rect 3074 11456 3126 11644
rect 3390 11456 3442 11644
rect -12146 9350 -11974 9726
rect -11786 9114 -11586 9962
rect -10740 9350 -10568 9726
rect -10380 9114 -10180 9962
rect -9334 9350 -9162 9726
rect -8974 9114 -8774 9962
rect -7928 9350 -7756 9726
rect -7568 9114 -7368 9962
rect 546 11146 598 11334
rect 862 11146 914 11334
rect 1178 11146 1230 11334
rect 1494 11146 1546 11334
rect 1810 11146 1862 11334
rect 2126 11146 2178 11334
rect 2442 11146 2494 11334
rect 2758 11146 2810 11334
rect 3074 11146 3126 11334
rect 3390 11146 3442 11334
rect 546 10838 598 11026
rect 862 10838 914 11026
rect 1178 10838 1230 11026
rect 1494 10838 1546 11026
rect 1810 10838 1862 11026
rect 2126 10838 2178 11026
rect 2442 10838 2494 11026
rect 2758 10838 2810 11026
rect 3074 10838 3126 11026
rect 3390 10838 3442 11026
rect 546 10526 598 10712
rect 862 10526 914 10712
rect 1178 10526 1230 10712
rect 1494 10526 1546 10712
rect 1810 10526 1862 10712
rect 2126 10526 2178 10712
rect 2442 10526 2494 10712
rect 2758 10526 2810 10712
rect 3074 10526 3126 10712
rect 3390 10526 3442 10712
rect 546 10218 598 10404
rect 862 10218 914 10404
rect 1178 10218 1230 10404
rect 1494 10218 1546 10404
rect 1810 10218 1862 10404
rect 2126 10218 2178 10404
rect 2442 10218 2494 10404
rect 2758 10218 2810 10404
rect 3074 10218 3126 10404
rect 3390 10218 3442 10404
rect 544 10038 3446 10046
rect 544 10002 3446 10038
rect 544 9994 3446 10002
rect -4168 8912 -3986 9236
rect -12146 7744 -11974 8120
rect -11786 7508 -11586 8356
rect -10740 7744 -10568 8120
rect -10380 7508 -10180 8356
rect -9334 7744 -9162 8120
rect -8974 7508 -8774 8356
rect -7928 7744 -7756 8120
rect -7568 7508 -7368 8356
rect -12146 6138 -11974 6514
rect -11786 5902 -11586 6750
rect -10740 6138 -10568 6514
rect -10380 5902 -10180 6750
rect -9334 6138 -9162 6514
rect -8974 5902 -8774 6750
rect -7928 6138 -7756 6514
rect -7568 5902 -7368 6750
<< metal2 >>
rect -1254 31608 9582 31618
rect -1254 31028 -1244 31608
rect 8992 31028 9582 31608
rect -1254 31018 9582 31028
rect -1254 30864 -654 31018
rect -454 30864 146 31018
rect 346 30864 946 31018
rect 1146 30864 1746 31018
rect 1946 30864 2546 31018
rect 2746 30864 3346 31018
rect 3546 30864 4146 31018
rect 4346 30864 7584 31018
rect -1532 30854 7584 30864
rect -1532 30274 -1522 30854
rect 7242 30274 7584 30854
rect -1532 30264 7584 30274
rect 3928 30186 4298 30264
rect 4586 30186 5186 30264
rect -1234 30080 -434 30090
rect -2992 30034 -2386 30044
rect -17432 29690 -3280 29700
rect -17432 29110 -17422 29690
rect -16842 29110 -16222 29690
rect -15642 29110 -15022 29690
rect -14442 29110 -13822 29690
rect -13242 29110 -12622 29690
rect -12042 29110 -11422 29690
rect -10842 29110 -10222 29690
rect -9642 29110 -9022 29690
rect -8442 29110 -7822 29690
rect -7242 29110 -6622 29690
rect -6042 29110 -5422 29690
rect -4842 29110 -3870 29690
rect -17432 29100 -3870 29110
rect -17430 29096 -17206 29100
rect -18166 28902 -17566 28910
rect -18166 27960 -18156 28902
rect -17580 27960 -17566 28902
rect -18166 27576 -17566 27960
rect -18166 26554 -18156 27576
rect -17580 26554 -17566 27576
rect -18166 26170 -17566 26554
rect -18166 25148 -18156 26170
rect -17580 25148 -17566 26170
rect -18166 24764 -17566 25148
rect -18166 23742 -18156 24764
rect -17580 23742 -17566 24764
rect -18166 23654 -17786 23742
rect -17590 23654 -17566 23742
rect -18166 23358 -17566 23654
rect -18166 22336 -18156 23358
rect -17580 22336 -17566 23358
rect -18166 22048 -17786 22336
rect -17590 22048 -17566 22336
rect -18166 21952 -17566 22048
rect -18166 20930 -18156 21952
rect -17580 20930 -17566 21952
rect -18166 20842 -17566 20930
rect -18166 20546 -17786 20842
rect -17590 20546 -17566 20842
rect -18166 19524 -18156 20546
rect -17580 19524 -17566 20546
rect -18166 19236 -17566 19524
rect -18166 19140 -17786 19236
rect -17590 19140 -17566 19236
rect -18166 18118 -18156 19140
rect -17580 18118 -17566 19140
rect -18166 17734 -17566 18118
rect -18166 16712 -18156 17734
rect -17580 16712 -17566 17734
rect -18166 16328 -17566 16712
rect -18166 15306 -18156 16328
rect -17580 15306 -17566 16328
rect -18166 14922 -17566 15306
rect -18166 13900 -18156 14922
rect -17580 13900 -17566 14922
rect -18166 13215 -17566 13900
rect -17430 28254 -17404 29096
rect -17222 28254 -17206 29096
rect -16024 29096 -15800 29100
rect -17430 27490 -17206 28254
rect -17430 26648 -17404 27490
rect -17222 26648 -17206 27490
rect -17430 25884 -17206 26648
rect -17430 25042 -17404 25884
rect -17222 25042 -17206 25884
rect -17430 24278 -17206 25042
rect -17430 23436 -17404 24278
rect -17222 23436 -17206 24278
rect -17430 22672 -17206 23436
rect -17430 21830 -17404 22672
rect -17222 21830 -17206 22672
rect -17430 21066 -17206 21830
rect -17430 20224 -17404 21066
rect -17222 20224 -17206 21066
rect -17430 19460 -17206 20224
rect -17430 18618 -17404 19460
rect -17222 18618 -17206 19460
rect -17430 17854 -17206 18618
rect -17430 17012 -17404 17854
rect -17222 17012 -17206 17854
rect -17430 16248 -17206 17012
rect -17430 15406 -17404 16248
rect -17222 15406 -17206 16248
rect -17430 14642 -17206 15406
rect -17430 13800 -17404 14642
rect -17222 13898 -17206 14642
rect -16760 28902 -16160 28910
rect -16760 27960 -16750 28902
rect -16174 27960 -16160 28902
rect -16760 27576 -16160 27960
rect -16760 26554 -16750 27576
rect -16174 26554 -16160 27576
rect -16760 26170 -16160 26554
rect -16760 25148 -16750 26170
rect -16174 25148 -16160 26170
rect -16760 24764 -16160 25148
rect -16760 23742 -16750 24764
rect -16174 23742 -16160 24764
rect -16760 23654 -16380 23742
rect -16184 23654 -16160 23742
rect -16760 23358 -16160 23654
rect -16760 22336 -16750 23358
rect -16174 22336 -16160 23358
rect -16760 22048 -16380 22336
rect -16184 22048 -16160 22336
rect -16760 21952 -16160 22048
rect -16760 20930 -16750 21952
rect -16174 20930 -16160 21952
rect -16760 20842 -16160 20930
rect -16760 20546 -16380 20842
rect -16184 20546 -16160 20842
rect -16760 19524 -16750 20546
rect -16174 19524 -16160 20546
rect -16760 19236 -16160 19524
rect -16760 19140 -16380 19236
rect -16184 19140 -16160 19236
rect -16760 18118 -16750 19140
rect -16174 18118 -16160 19140
rect -16760 17734 -16160 18118
rect -16760 16712 -16750 17734
rect -16174 16712 -16160 17734
rect -16760 16328 -16160 16712
rect -16760 15306 -16750 16328
rect -16174 15306 -16160 16328
rect -16760 14922 -16160 15306
rect -16760 13900 -16750 14922
rect -16174 13900 -16160 14922
rect -17222 13800 -17208 13898
rect -17430 13594 -17208 13800
rect -18166 13212 -17226 13215
rect -16760 13212 -16160 13900
rect -16024 28254 -15998 29096
rect -15816 28254 -15800 29096
rect -14618 29096 -14394 29100
rect -16024 27490 -15800 28254
rect -16024 26648 -15998 27490
rect -15816 26648 -15800 27490
rect -16024 25884 -15800 26648
rect -16024 25042 -15998 25884
rect -15816 25042 -15800 25884
rect -16024 24278 -15800 25042
rect -16024 23436 -15998 24278
rect -15816 23436 -15800 24278
rect -16024 22672 -15800 23436
rect -16024 21830 -15998 22672
rect -15816 21830 -15800 22672
rect -16024 21066 -15800 21830
rect -16024 20224 -15998 21066
rect -15816 20224 -15800 21066
rect -16024 19460 -15800 20224
rect -16024 18618 -15998 19460
rect -15816 18618 -15800 19460
rect -16024 17854 -15800 18618
rect -16024 17012 -15998 17854
rect -15816 17012 -15800 17854
rect -16024 16248 -15800 17012
rect -16024 15406 -15998 16248
rect -15816 15406 -15800 16248
rect -16024 14642 -15800 15406
rect -16024 13800 -15998 14642
rect -15816 13898 -15800 14642
rect -15354 28902 -14754 28910
rect -15354 27960 -15344 28902
rect -14768 27960 -14754 28902
rect -15354 27576 -14754 27960
rect -15354 26554 -15344 27576
rect -14768 26554 -14754 27576
rect -15354 26170 -14754 26554
rect -15354 25148 -15344 26170
rect -14768 25148 -14754 26170
rect -15354 24764 -14754 25148
rect -15354 23742 -15344 24764
rect -14768 23742 -14754 24764
rect -15354 23654 -14974 23742
rect -14778 23654 -14754 23742
rect -15354 23358 -14754 23654
rect -15354 22336 -15344 23358
rect -14768 22336 -14754 23358
rect -15354 22048 -14974 22336
rect -14778 22048 -14754 22336
rect -15354 21952 -14754 22048
rect -15354 20930 -15344 21952
rect -14768 20930 -14754 21952
rect -15354 20842 -14754 20930
rect -15354 20546 -14974 20842
rect -14778 20546 -14754 20842
rect -15354 19524 -15344 20546
rect -14768 19524 -14754 20546
rect -15354 19236 -14754 19524
rect -15354 19140 -14974 19236
rect -14778 19140 -14754 19236
rect -15354 18118 -15344 19140
rect -14768 18118 -14754 19140
rect -15354 17734 -14754 18118
rect -15354 16712 -15344 17734
rect -14768 16712 -14754 17734
rect -15354 16328 -14754 16712
rect -15354 15306 -15344 16328
rect -14768 15306 -14754 16328
rect -15354 14922 -14754 15306
rect -15354 13900 -15344 14922
rect -14768 13900 -14754 14922
rect -15816 13800 -15802 13898
rect -16024 13594 -15802 13800
rect -15354 13212 -14754 13900
rect -14618 28254 -14592 29096
rect -14410 28254 -14394 29096
rect -13212 29096 -12988 29100
rect -14618 27490 -14394 28254
rect -14618 26648 -14592 27490
rect -14410 26648 -14394 27490
rect -14618 25884 -14394 26648
rect -14618 25042 -14592 25884
rect -14410 25042 -14394 25884
rect -14618 24278 -14394 25042
rect -14618 23436 -14592 24278
rect -14410 23436 -14394 24278
rect -14618 22672 -14394 23436
rect -14618 21830 -14592 22672
rect -14410 21830 -14394 22672
rect -14618 21066 -14394 21830
rect -14618 20224 -14592 21066
rect -14410 20224 -14394 21066
rect -14618 19460 -14394 20224
rect -14618 18618 -14592 19460
rect -14410 18618 -14394 19460
rect -14618 17854 -14394 18618
rect -14618 17012 -14592 17854
rect -14410 17012 -14394 17854
rect -14618 16248 -14394 17012
rect -14618 15406 -14592 16248
rect -14410 15406 -14394 16248
rect -14618 14642 -14394 15406
rect -14618 13800 -14592 14642
rect -14410 13898 -14394 14642
rect -13948 28902 -13348 28910
rect -13948 27960 -13938 28902
rect -13362 27960 -13348 28902
rect -13948 27576 -13348 27960
rect -13948 26554 -13938 27576
rect -13362 26554 -13348 27576
rect -13948 26170 -13348 26554
rect -13948 25148 -13938 26170
rect -13362 25148 -13348 26170
rect -13948 24764 -13348 25148
rect -13948 23742 -13938 24764
rect -13362 23742 -13348 24764
rect -13948 23654 -13568 23742
rect -13372 23654 -13348 23742
rect -13948 23358 -13348 23654
rect -13948 22336 -13938 23358
rect -13362 22336 -13348 23358
rect -13948 22048 -13568 22336
rect -13372 22048 -13348 22336
rect -13948 21952 -13348 22048
rect -13948 20930 -13938 21952
rect -13362 20930 -13348 21952
rect -13948 20842 -13348 20930
rect -13948 20546 -13568 20842
rect -13372 20546 -13348 20842
rect -13948 19524 -13938 20546
rect -13362 19524 -13348 20546
rect -13948 19236 -13348 19524
rect -13948 19140 -13568 19236
rect -13372 19140 -13348 19236
rect -13948 18118 -13938 19140
rect -13362 18118 -13348 19140
rect -13948 17734 -13348 18118
rect -13948 16712 -13938 17734
rect -13362 16712 -13348 17734
rect -13948 16328 -13348 16712
rect -13948 15306 -13938 16328
rect -13362 15306 -13348 16328
rect -13948 14922 -13348 15306
rect -13948 13900 -13938 14922
rect -13362 13900 -13348 14922
rect -14410 13800 -14396 13898
rect -14618 13594 -14396 13800
rect -13948 13212 -13348 13900
rect -13212 28254 -13186 29096
rect -13004 28254 -12988 29096
rect -11806 29096 -11582 29100
rect -13212 27490 -12988 28254
rect -13212 26648 -13186 27490
rect -13004 26648 -12988 27490
rect -13212 25884 -12988 26648
rect -13212 25042 -13186 25884
rect -13004 25042 -12988 25884
rect -13212 24278 -12988 25042
rect -13212 23436 -13186 24278
rect -13004 23436 -12988 24278
rect -13212 22672 -12988 23436
rect -13212 21830 -13186 22672
rect -13004 21830 -12988 22672
rect -13212 21066 -12988 21830
rect -13212 20224 -13186 21066
rect -13004 20224 -12988 21066
rect -13212 19460 -12988 20224
rect -13212 18618 -13186 19460
rect -13004 18618 -12988 19460
rect -13212 17854 -12988 18618
rect -13212 17012 -13186 17854
rect -13004 17012 -12988 17854
rect -13212 16248 -12988 17012
rect -13212 15406 -13186 16248
rect -13004 15406 -12988 16248
rect -13212 14642 -12988 15406
rect -13212 13800 -13186 14642
rect -13004 13898 -12988 14642
rect -12542 28902 -11942 28910
rect -12542 27960 -12532 28902
rect -11956 27960 -11942 28902
rect -12542 27576 -11942 27960
rect -12542 26554 -12532 27576
rect -11956 26554 -11942 27576
rect -12542 26170 -11942 26554
rect -12542 25148 -12532 26170
rect -11956 25148 -11942 26170
rect -12542 24764 -11942 25148
rect -12542 23742 -12532 24764
rect -11956 23742 -11942 24764
rect -12542 23654 -12162 23742
rect -11966 23654 -11942 23742
rect -12542 23358 -11942 23654
rect -12542 22336 -12532 23358
rect -11956 22336 -11942 23358
rect -12542 22048 -12162 22336
rect -11966 22048 -11942 22336
rect -12542 21952 -11942 22048
rect -12542 20930 -12532 21952
rect -11956 20930 -11942 21952
rect -12542 20842 -11942 20930
rect -12542 20546 -12162 20842
rect -11966 20546 -11942 20842
rect -12542 19524 -12532 20546
rect -11956 19524 -11942 20546
rect -12542 19236 -11942 19524
rect -12542 19140 -12162 19236
rect -11966 19140 -11942 19236
rect -12542 18118 -12532 19140
rect -11956 18118 -11942 19140
rect -12542 17734 -11942 18118
rect -12542 16712 -12532 17734
rect -11956 16712 -11942 17734
rect -12542 16328 -11942 16712
rect -12542 15306 -12532 16328
rect -11956 15306 -11942 16328
rect -12542 14922 -11942 15306
rect -12542 13900 -12532 14922
rect -11956 13900 -11942 14922
rect -13004 13800 -12990 13898
rect -13212 13594 -12990 13800
rect -12542 13212 -11942 13900
rect -11806 28254 -11780 29096
rect -11598 28254 -11582 29096
rect -10400 29096 -10176 29100
rect -11806 27490 -11582 28254
rect -11806 26648 -11780 27490
rect -11598 26648 -11582 27490
rect -11806 25884 -11582 26648
rect -11806 25042 -11780 25884
rect -11598 25042 -11582 25884
rect -11806 24278 -11582 25042
rect -11806 23436 -11780 24278
rect -11598 23436 -11582 24278
rect -11806 22672 -11582 23436
rect -11806 21830 -11780 22672
rect -11598 21830 -11582 22672
rect -11806 21066 -11582 21830
rect -11806 20224 -11780 21066
rect -11598 20224 -11582 21066
rect -11806 19460 -11582 20224
rect -11806 18618 -11780 19460
rect -11598 18618 -11582 19460
rect -11806 17854 -11582 18618
rect -11806 17012 -11780 17854
rect -11598 17012 -11582 17854
rect -11806 16248 -11582 17012
rect -11806 15406 -11780 16248
rect -11598 15406 -11582 16248
rect -11806 14642 -11582 15406
rect -11806 13800 -11780 14642
rect -11598 13898 -11582 14642
rect -11136 28902 -10536 28910
rect -11136 27960 -11126 28902
rect -10550 27960 -10536 28902
rect -11136 27576 -10536 27960
rect -11136 26554 -11126 27576
rect -10550 26554 -10536 27576
rect -11136 26170 -10536 26554
rect -11136 25148 -11126 26170
rect -10550 25148 -10536 26170
rect -11136 24764 -10536 25148
rect -11136 23742 -11126 24764
rect -10550 23742 -10536 24764
rect -11136 23654 -10756 23742
rect -10560 23654 -10536 23742
rect -11136 23358 -10536 23654
rect -11136 22336 -11126 23358
rect -10550 22336 -10536 23358
rect -11136 22048 -10756 22336
rect -10560 22048 -10536 22336
rect -11136 21952 -10536 22048
rect -11136 20930 -11126 21952
rect -10550 20930 -10536 21952
rect -11136 20842 -10536 20930
rect -11136 20546 -10756 20842
rect -10560 20546 -10536 20842
rect -11136 19524 -11126 20546
rect -10550 19524 -10536 20546
rect -11136 19236 -10536 19524
rect -11136 19140 -10756 19236
rect -10560 19140 -10536 19236
rect -11136 18118 -11126 19140
rect -10550 18118 -10536 19140
rect -11136 17734 -10536 18118
rect -11136 16712 -11126 17734
rect -10550 16712 -10536 17734
rect -11136 16328 -10536 16712
rect -11136 15306 -11126 16328
rect -10550 15306 -10536 16328
rect -11136 14922 -10536 15306
rect -11136 13900 -11126 14922
rect -10550 13900 -10536 14922
rect -11598 13800 -11584 13898
rect -11806 13594 -11584 13800
rect -11136 13212 -10536 13900
rect -10400 28254 -10374 29096
rect -10192 28254 -10176 29096
rect -8994 29096 -8770 29100
rect -10400 27490 -10176 28254
rect -10400 26648 -10374 27490
rect -10192 26648 -10176 27490
rect -10400 25884 -10176 26648
rect -10400 25042 -10374 25884
rect -10192 25042 -10176 25884
rect -10400 24278 -10176 25042
rect -10400 23436 -10374 24278
rect -10192 23436 -10176 24278
rect -10400 22672 -10176 23436
rect -10400 21830 -10374 22672
rect -10192 21830 -10176 22672
rect -10400 21066 -10176 21830
rect -10400 20224 -10374 21066
rect -10192 20224 -10176 21066
rect -10400 19460 -10176 20224
rect -10400 18618 -10374 19460
rect -10192 18618 -10176 19460
rect -10400 17854 -10176 18618
rect -10400 17012 -10374 17854
rect -10192 17012 -10176 17854
rect -10400 16248 -10176 17012
rect -10400 15406 -10374 16248
rect -10192 15406 -10176 16248
rect -10400 14642 -10176 15406
rect -10400 13800 -10374 14642
rect -10192 13898 -10176 14642
rect -9730 28902 -9130 28910
rect -9730 27960 -9720 28902
rect -9144 27960 -9130 28902
rect -9730 27576 -9130 27960
rect -9730 26554 -9720 27576
rect -9144 26554 -9130 27576
rect -9730 26170 -9130 26554
rect -9730 25148 -9720 26170
rect -9144 25148 -9130 26170
rect -9730 24764 -9130 25148
rect -9730 23742 -9720 24764
rect -9144 23742 -9130 24764
rect -9730 23654 -9350 23742
rect -9154 23654 -9130 23742
rect -9730 23358 -9130 23654
rect -9730 22336 -9720 23358
rect -9144 22336 -9130 23358
rect -9730 22048 -9350 22336
rect -9154 22048 -9130 22336
rect -9730 21952 -9130 22048
rect -9730 20930 -9720 21952
rect -9144 20930 -9130 21952
rect -9730 20842 -9130 20930
rect -9730 20546 -9350 20842
rect -9154 20546 -9130 20842
rect -9730 19524 -9720 20546
rect -9144 19524 -9130 20546
rect -9730 19236 -9130 19524
rect -9730 19140 -9350 19236
rect -9154 19140 -9130 19236
rect -9730 18118 -9720 19140
rect -9144 18118 -9130 19140
rect -9730 17734 -9130 18118
rect -9730 16712 -9720 17734
rect -9144 16712 -9130 17734
rect -9730 16328 -9130 16712
rect -9730 15306 -9720 16328
rect -9144 15306 -9130 16328
rect -9730 14922 -9130 15306
rect -9730 13900 -9720 14922
rect -9144 13900 -9130 14922
rect -10192 13800 -10178 13898
rect -10400 13594 -10178 13800
rect -9730 13212 -9130 13900
rect -8994 28254 -8968 29096
rect -8786 28254 -8770 29096
rect -7588 29096 -7364 29100
rect -8994 27490 -8770 28254
rect -8994 26648 -8968 27490
rect -8786 26648 -8770 27490
rect -8994 25884 -8770 26648
rect -8994 25042 -8968 25884
rect -8786 25042 -8770 25884
rect -8994 24278 -8770 25042
rect -8994 23436 -8968 24278
rect -8786 23436 -8770 24278
rect -8994 22672 -8770 23436
rect -8994 21830 -8968 22672
rect -8786 21830 -8770 22672
rect -8994 21066 -8770 21830
rect -8994 20224 -8968 21066
rect -8786 20224 -8770 21066
rect -8994 19460 -8770 20224
rect -8994 18618 -8968 19460
rect -8786 18618 -8770 19460
rect -8994 17854 -8770 18618
rect -8994 17012 -8968 17854
rect -8786 17012 -8770 17854
rect -8994 16248 -8770 17012
rect -8994 15406 -8968 16248
rect -8786 15406 -8770 16248
rect -8994 14642 -8770 15406
rect -8994 13800 -8968 14642
rect -8786 13898 -8770 14642
rect -8324 28902 -7724 28910
rect -8324 27960 -8314 28902
rect -7738 27960 -7724 28902
rect -8324 27576 -7724 27960
rect -8324 26554 -8314 27576
rect -7738 26554 -7724 27576
rect -8324 26170 -7724 26554
rect -8324 25148 -8314 26170
rect -7738 25148 -7724 26170
rect -8324 24764 -7724 25148
rect -8324 23742 -8314 24764
rect -7738 23742 -7724 24764
rect -8324 23654 -7944 23742
rect -7748 23654 -7724 23742
rect -8324 23358 -7724 23654
rect -8324 22336 -8314 23358
rect -7738 22336 -7724 23358
rect -8324 22048 -7944 22336
rect -7748 22048 -7724 22336
rect -8324 21952 -7724 22048
rect -8324 20930 -8314 21952
rect -7738 20930 -7724 21952
rect -8324 20842 -7724 20930
rect -8324 20546 -7944 20842
rect -7748 20546 -7724 20842
rect -8324 19524 -8314 20546
rect -7738 19524 -7724 20546
rect -8324 19236 -7724 19524
rect -8324 19140 -7944 19236
rect -7748 19140 -7724 19236
rect -8324 18118 -8314 19140
rect -7738 18118 -7724 19140
rect -8324 17734 -7724 18118
rect -8324 16712 -8314 17734
rect -7738 16712 -7724 17734
rect -8324 16328 -7724 16712
rect -8324 15306 -8314 16328
rect -7738 15306 -7724 16328
rect -8324 14922 -7724 15306
rect -8324 13900 -8314 14922
rect -7738 13900 -7724 14922
rect -8786 13800 -8772 13898
rect -8994 13594 -8772 13800
rect -8324 13212 -7724 13900
rect -7588 28254 -7562 29096
rect -7380 28254 -7364 29096
rect -6182 29096 -5958 29100
rect -7588 27490 -7364 28254
rect -7588 26648 -7562 27490
rect -7380 26648 -7364 27490
rect -7588 25884 -7364 26648
rect -7588 25042 -7562 25884
rect -7380 25042 -7364 25884
rect -7588 24278 -7364 25042
rect -7588 23436 -7562 24278
rect -7380 23436 -7364 24278
rect -7588 22672 -7364 23436
rect -7588 21830 -7562 22672
rect -7380 21830 -7364 22672
rect -7588 21066 -7364 21830
rect -7588 20224 -7562 21066
rect -7380 20224 -7364 21066
rect -7588 19460 -7364 20224
rect -7588 18618 -7562 19460
rect -7380 18618 -7364 19460
rect -7588 17854 -7364 18618
rect -7588 17012 -7562 17854
rect -7380 17012 -7364 17854
rect -7588 16248 -7364 17012
rect -7588 15406 -7562 16248
rect -7380 15406 -7364 16248
rect -7588 14642 -7364 15406
rect -7588 13800 -7562 14642
rect -7380 13898 -7364 14642
rect -6918 28902 -6318 28910
rect -6918 27960 -6908 28902
rect -6332 27960 -6318 28902
rect -6918 27576 -6318 27960
rect -6918 26554 -6908 27576
rect -6332 26554 -6318 27576
rect -6918 26170 -6318 26554
rect -6918 25148 -6908 26170
rect -6332 25148 -6318 26170
rect -6918 24764 -6318 25148
rect -6918 23742 -6908 24764
rect -6332 23742 -6318 24764
rect -6918 23654 -6538 23742
rect -6342 23654 -6318 23742
rect -6918 23358 -6318 23654
rect -6918 22336 -6908 23358
rect -6332 22336 -6318 23358
rect -6918 22048 -6538 22336
rect -6342 22048 -6318 22336
rect -6918 21952 -6318 22048
rect -6918 20930 -6908 21952
rect -6332 20930 -6318 21952
rect -6918 20842 -6318 20930
rect -6918 20546 -6538 20842
rect -6342 20546 -6318 20842
rect -6918 19524 -6908 20546
rect -6332 19524 -6318 20546
rect -6918 19236 -6318 19524
rect -6918 19140 -6538 19236
rect -6342 19140 -6318 19236
rect -6918 18118 -6908 19140
rect -6332 18118 -6318 19140
rect -6918 17734 -6318 18118
rect -6918 16712 -6908 17734
rect -6332 16712 -6318 17734
rect -6918 16328 -6318 16712
rect -6918 15306 -6908 16328
rect -6332 15306 -6318 16328
rect -6918 14922 -6318 15306
rect -6918 13900 -6908 14922
rect -6332 13900 -6318 14922
rect -7380 13800 -7366 13898
rect -7588 13594 -7366 13800
rect -6918 13212 -6318 13900
rect -6182 28254 -6156 29096
rect -5974 28254 -5958 29096
rect -4776 29096 -4552 29100
rect -6182 27490 -5958 28254
rect -6182 26648 -6156 27490
rect -5974 26648 -5958 27490
rect -6182 25884 -5958 26648
rect -6182 25042 -6156 25884
rect -5974 25042 -5958 25884
rect -6182 24278 -5958 25042
rect -6182 23436 -6156 24278
rect -5974 23436 -5958 24278
rect -6182 22672 -5958 23436
rect -6182 21830 -6156 22672
rect -5974 21830 -5958 22672
rect -6182 21066 -5958 21830
rect -6182 20224 -6156 21066
rect -5974 20224 -5958 21066
rect -6182 19460 -5958 20224
rect -6182 18618 -6156 19460
rect -5974 18618 -5958 19460
rect -6182 17854 -5958 18618
rect -6182 17012 -6156 17854
rect -5974 17012 -5958 17854
rect -6182 16248 -5958 17012
rect -6182 15406 -6156 16248
rect -5974 15406 -5958 16248
rect -6182 14642 -5958 15406
rect -6182 13800 -6156 14642
rect -5974 13898 -5958 14642
rect -5512 28902 -4912 28910
rect -5512 27960 -5502 28902
rect -4926 27960 -4912 28902
rect -5512 27576 -4912 27960
rect -5512 26554 -5502 27576
rect -4926 26554 -4912 27576
rect -5512 26170 -4912 26554
rect -5512 25148 -5502 26170
rect -4926 25148 -4912 26170
rect -5512 24764 -4912 25148
rect -5512 23742 -5502 24764
rect -4926 23742 -4912 24764
rect -5512 23654 -5132 23742
rect -4936 23654 -4912 23742
rect -5512 23358 -4912 23654
rect -5512 22336 -5502 23358
rect -4926 22336 -4912 23358
rect -5512 22048 -5132 22336
rect -4936 22048 -4912 22336
rect -5512 21952 -4912 22048
rect -5512 20930 -5502 21952
rect -4926 20930 -4912 21952
rect -5512 20842 -4912 20930
rect -5512 20546 -5132 20842
rect -4936 20546 -4912 20842
rect -5512 19524 -5502 20546
rect -4926 19524 -4912 20546
rect -5512 19236 -4912 19524
rect -5512 19140 -5132 19236
rect -4936 19140 -4912 19236
rect -5512 18118 -5502 19140
rect -4926 18118 -4912 19140
rect -5512 17734 -4912 18118
rect -5512 16712 -5502 17734
rect -4926 16712 -4912 17734
rect -5512 16328 -4912 16712
rect -5512 15306 -5502 16328
rect -4926 15306 -4912 16328
rect -5512 14922 -4912 15306
rect -5512 13900 -5502 14922
rect -4926 13900 -4912 14922
rect -5974 13800 -5960 13898
rect -6182 13594 -5960 13800
rect -5512 13212 -4912 13900
rect -4776 28254 -4750 29096
rect -4568 28254 -4552 29096
rect -4776 27490 -4552 28254
rect -4776 26648 -4750 27490
rect -4568 26648 -4552 27490
rect -4776 25884 -4552 26648
rect -4776 25042 -4750 25884
rect -4568 25042 -4552 25884
rect -4776 24278 -4552 25042
rect -4776 23436 -4750 24278
rect -4568 23436 -4552 24278
rect -4776 22672 -4552 23436
rect -4776 21830 -4750 22672
rect -4568 21830 -4552 22672
rect -4776 21066 -4552 21830
rect -4776 20224 -4750 21066
rect -4568 20224 -4552 21066
rect -4776 19460 -4552 20224
rect -4776 18618 -4750 19460
rect -4568 18618 -4552 19460
rect -4776 17854 -4552 18618
rect -4776 17012 -4750 17854
rect -4568 17012 -4552 17854
rect -4776 16248 -4552 17012
rect -4776 15406 -4750 16248
rect -4568 15406 -4552 16248
rect -4776 14642 -4552 15406
rect -4776 13800 -4750 14642
rect -4568 13800 -4552 14642
rect -4776 13594 -4552 13800
rect -3880 28490 -3870 29100
rect -3290 28490 -3280 29690
rect -18166 13206 -4912 13212
rect -18166 13202 -17826 13206
rect -17226 13202 -16826 13206
rect -16160 13202 -15826 13206
rect -14226 13202 -13948 13206
rect -13226 13202 -12826 13206
rect -11942 13202 -11826 13206
rect -11226 13202 -11136 13206
rect -10226 13202 -9826 13206
rect -9130 13202 -8826 13206
rect -7226 13202 -6918 13206
rect -6226 13202 -5826 13206
rect -18166 12606 -18156 13202
rect -18166 12596 -4912 12606
rect -3880 12886 -3280 28490
rect -2992 24656 -2982 30034
rect -2396 29990 -2386 30034
rect -1234 29990 -1224 30080
rect -2396 29390 -1224 29990
rect -2396 28594 -2386 29390
rect -1234 29300 -1224 29390
rect -444 29990 -434 30080
rect 162 30080 962 30090
rect 162 29990 172 30080
rect -444 29390 172 29990
rect -444 29300 -434 29390
rect -1234 29290 -434 29300
rect 162 29300 172 29390
rect 952 29990 962 30080
rect 1558 30080 2358 30090
rect 1558 29990 1568 30080
rect 952 29390 1568 29990
rect 952 29300 962 29390
rect 162 29290 962 29300
rect 1558 29300 1568 29390
rect 2348 29990 2358 30080
rect 2954 30080 3754 30090
rect 2954 29990 2964 30080
rect 2348 29390 2964 29990
rect 2348 29300 2358 29390
rect 1558 29290 2358 29300
rect 2954 29300 2964 29390
rect 3744 29300 3754 30080
rect 2954 29290 3754 29300
rect 3928 29586 5186 30186
rect 3928 29386 4298 29586
rect 5384 29386 5984 30264
rect 3928 29116 5984 29386
rect -1780 29106 5984 29116
rect -1780 28878 -1696 29106
rect -1368 28878 -300 29106
rect 28 28878 1096 29106
rect 1424 28878 2492 29106
rect 2820 28878 3888 29106
rect 4216 28878 5984 29106
rect -1780 28868 5984 28878
rect 3928 28786 5984 28868
rect -1234 28684 -434 28694
rect -1234 28594 -1224 28684
rect -2396 27994 -1224 28594
rect -2396 27198 -2386 27994
rect -1234 27904 -1224 27994
rect -444 28594 -434 28684
rect 162 28684 962 28694
rect 162 28594 172 28684
rect -444 27994 172 28594
rect -444 27904 -434 27994
rect -1234 27894 -434 27904
rect 162 27904 172 27994
rect 952 28594 962 28684
rect 1558 28684 2358 28694
rect 1558 28594 1568 28684
rect 952 27994 1568 28594
rect 952 27904 962 27994
rect 162 27894 962 27904
rect 1558 27904 1568 27994
rect 2348 28594 2358 28684
rect 2954 28684 3754 28694
rect 2954 28594 2964 28684
rect 2348 27994 2964 28594
rect 2348 27904 2358 27994
rect 1558 27894 2358 27904
rect 2954 27904 2964 27994
rect 3744 27904 3754 28684
rect 2954 27894 3754 27904
rect 3928 28586 4298 28786
rect 5384 28784 5984 28786
rect 6184 28586 6784 30264
rect 3928 27986 6784 28586
rect 3928 27786 4298 27986
rect 6184 27984 6784 27986
rect 6984 27786 7584 30264
rect 3928 27720 7584 27786
rect -1780 27710 7584 27720
rect -1780 27482 -1696 27710
rect -1368 27482 -300 27710
rect 28 27482 1096 27710
rect 1424 27482 2492 27710
rect 2820 27482 3888 27710
rect 4216 27482 7584 27710
rect -1780 27472 7584 27482
rect -1234 27288 -434 27298
rect -1234 27198 -1224 27288
rect -2396 26598 -1224 27198
rect -2396 25802 -2386 26598
rect -1234 26508 -1224 26598
rect -444 27198 -434 27288
rect 162 27288 962 27298
rect 162 27198 172 27288
rect -444 26598 172 27198
rect -444 26508 -434 26598
rect -1234 26498 -434 26508
rect 162 26508 172 26598
rect 952 27198 962 27288
rect 1558 27288 2358 27298
rect 1558 27198 1568 27288
rect 952 26598 1568 27198
rect 952 26508 962 26598
rect 162 26498 962 26508
rect 1558 26508 1568 26598
rect 2348 27198 2358 27288
rect 2954 27288 3754 27298
rect 2954 27198 2964 27288
rect 2348 26598 2964 27198
rect 2348 26508 2358 26598
rect 1558 26498 2358 26508
rect 2954 26508 2964 26598
rect 3744 26508 3754 27288
rect 2954 26498 3754 26508
rect 3928 27186 7584 27472
rect 3928 26986 4298 27186
rect 6984 27184 7584 27186
rect 7784 26986 8384 31018
rect 8982 29318 9582 31018
rect 8982 29308 50192 29318
rect 8982 28728 8992 29308
rect 50182 28728 50192 29308
rect 8982 28718 50192 28728
rect 10784 28256 11032 28718
rect 9910 28166 10510 28200
rect 9910 28132 9920 28166
rect 9810 28122 9920 28132
rect 10500 28132 10510 28166
rect 10500 28122 10610 28132
rect 9810 27342 9820 28122
rect 10600 27342 10610 28122
rect 9810 27332 9920 27342
rect 3928 26386 8384 26986
rect 9910 26736 9920 27332
rect 3928 26324 4298 26386
rect 7784 26384 8384 26386
rect 9810 26726 9920 26736
rect 10500 27332 10610 27342
rect 10500 26736 10510 27332
rect 10500 26726 10610 26736
rect -1780 26314 4298 26324
rect -1780 26086 -1696 26314
rect -1368 26086 -300 26314
rect 28 26086 1096 26314
rect 1424 26086 2492 26314
rect 2820 26086 3888 26314
rect 4216 26086 4298 26314
rect -1780 26076 4298 26086
rect -1234 25892 -434 25902
rect -1234 25802 -1224 25892
rect -2396 25202 -1224 25802
rect -2396 24656 -2386 25202
rect -1234 25112 -1224 25202
rect -444 25802 -434 25892
rect 162 25892 962 25902
rect 162 25802 172 25892
rect -444 25202 172 25802
rect -444 25112 -434 25202
rect -1234 25102 -434 25112
rect 162 25112 172 25202
rect 952 25802 962 25892
rect 1558 25892 2358 25902
rect 1558 25802 1568 25892
rect 952 25202 1568 25802
rect 952 25112 962 25202
rect 162 25102 962 25112
rect 1558 25112 1568 25202
rect 2348 25802 2358 25892
rect 2954 25892 3754 25902
rect 2954 25802 2964 25892
rect 2348 25202 2964 25802
rect 2348 25112 2358 25202
rect 1558 25102 2358 25112
rect 2954 25112 2964 25202
rect 3744 25112 3754 25892
rect 2954 25102 3754 25112
rect 3928 24928 4298 26076
rect 9810 25946 9820 26726
rect 10600 25946 10610 26726
rect 9810 25936 9920 25946
rect -2992 24448 -2386 24656
rect -1780 24918 4298 24928
rect -1780 24690 -1696 24918
rect -1368 24690 -300 24918
rect 28 24690 1096 24918
rect 1424 24690 2492 24918
rect 2820 24690 3888 24918
rect 4216 24690 4298 24918
rect 9910 24784 9920 25936
rect -1780 24556 4298 24690
rect 4632 24774 9920 24784
rect 10500 25936 10610 25946
rect 10500 24784 10510 25936
rect 10784 25716 10796 28256
rect 11020 25716 11032 28256
rect 12180 28256 12428 28718
rect 11306 28166 11906 28200
rect 11306 28132 11316 28166
rect 11206 28122 11316 28132
rect 11896 28132 11906 28166
rect 11896 28122 12006 28132
rect 11206 27342 11216 28122
rect 11996 27342 12006 28122
rect 11206 27332 11316 27342
rect 11306 26736 11316 27332
rect 11206 26726 11316 26736
rect 11896 27332 12006 27342
rect 11896 26736 11906 27332
rect 11896 26726 12006 26736
rect 11206 25946 11216 26726
rect 11996 25946 12006 26726
rect 11206 25936 11316 25946
rect 10784 25704 11032 25716
rect 11306 24784 11316 25936
rect 10500 24774 11316 24784
rect 11896 25936 12006 25946
rect 11896 24784 11906 25936
rect 12180 25716 12192 28256
rect 12416 25716 12428 28256
rect 13576 28256 13824 28718
rect 12702 28166 13302 28200
rect 12702 28132 12712 28166
rect 12602 28122 12712 28132
rect 13292 28132 13302 28166
rect 13292 28122 13402 28132
rect 12602 27342 12612 28122
rect 13392 27342 13402 28122
rect 12602 27332 12712 27342
rect 12702 26736 12712 27332
rect 12602 26726 12712 26736
rect 13292 27332 13402 27342
rect 13292 26736 13302 27332
rect 13292 26726 13402 26736
rect 12602 25946 12612 26726
rect 13392 25946 13402 26726
rect 12602 25936 12712 25946
rect 12180 25704 12428 25716
rect 12702 24784 12712 25936
rect 11896 24774 12712 24784
rect 13292 25936 13402 25946
rect 13292 24784 13302 25936
rect 13576 25716 13588 28256
rect 13812 25716 13824 28256
rect 14972 28256 15220 28718
rect 14098 28166 14698 28200
rect 14098 28132 14108 28166
rect 13998 28122 14108 28132
rect 14688 28132 14698 28166
rect 14688 28122 14798 28132
rect 13998 27342 14008 28122
rect 14788 27342 14798 28122
rect 13998 27332 14108 27342
rect 14098 26736 14108 27332
rect 13998 26726 14108 26736
rect 14688 27332 14798 27342
rect 14688 26736 14698 27332
rect 14688 26726 14798 26736
rect 13998 25946 14008 26726
rect 14788 25946 14798 26726
rect 13998 25936 14108 25946
rect 13576 25704 13824 25716
rect 14098 24784 14108 25936
rect 13292 24774 14108 24784
rect 14688 25936 14798 25946
rect 14688 24784 14698 25936
rect 14972 25716 14984 28256
rect 15208 25716 15220 28256
rect 16368 28256 16616 28718
rect 15494 28166 16094 28200
rect 15494 28132 15504 28166
rect 15394 28122 15504 28132
rect 16084 28132 16094 28166
rect 16084 28122 16194 28132
rect 15394 27342 15404 28122
rect 16184 27342 16194 28122
rect 15394 27332 15504 27342
rect 15494 26736 15504 27332
rect 15394 26726 15504 26736
rect 16084 27332 16194 27342
rect 16084 26736 16094 27332
rect 16084 26726 16194 26736
rect 15394 25946 15404 26726
rect 16184 25946 16194 26726
rect 15394 25936 15504 25946
rect 14972 25704 15220 25716
rect 15494 24784 15504 25936
rect 14688 24774 15504 24784
rect 16084 25936 16194 25946
rect 16084 24784 16094 25936
rect 16368 25716 16380 28256
rect 16604 25716 16616 28256
rect 17764 28256 18012 28718
rect 16890 28166 17490 28200
rect 16890 28132 16900 28166
rect 16790 28122 16900 28132
rect 17480 28132 17490 28166
rect 17480 28122 17590 28132
rect 16790 27342 16800 28122
rect 17580 27342 17590 28122
rect 16790 27332 16900 27342
rect 16890 26736 16900 27332
rect 16790 26726 16900 26736
rect 17480 27332 17590 27342
rect 17480 26736 17490 27332
rect 17480 26726 17590 26736
rect 16790 25946 16800 26726
rect 17580 25946 17590 26726
rect 16790 25936 16900 25946
rect 16368 25704 16616 25716
rect 16890 24784 16900 25936
rect 16084 24774 16900 24784
rect 17480 25936 17590 25946
rect 17480 24784 17490 25936
rect 17764 25716 17776 28256
rect 18000 25716 18012 28256
rect 19160 28256 19408 28718
rect 18286 28166 18886 28200
rect 18286 28132 18296 28166
rect 18186 28122 18296 28132
rect 18876 28132 18886 28166
rect 18876 28122 18986 28132
rect 18186 27342 18196 28122
rect 18976 27342 18986 28122
rect 18186 27332 18296 27342
rect 18286 26736 18296 27332
rect 18186 26726 18296 26736
rect 18876 27332 18986 27342
rect 18876 26736 18886 27332
rect 18876 26726 18986 26736
rect 18186 25946 18196 26726
rect 18976 25946 18986 26726
rect 18186 25936 18296 25946
rect 17764 25704 18012 25716
rect 18286 24784 18296 25936
rect 17480 24774 18296 24784
rect 18876 25936 18986 25946
rect 18876 24784 18886 25936
rect 19160 25716 19172 28256
rect 19396 25716 19408 28256
rect 20556 28256 20804 28718
rect 19682 28166 20282 28200
rect 19682 28132 19692 28166
rect 19582 28122 19692 28132
rect 20272 28132 20282 28166
rect 20272 28122 20382 28132
rect 19582 27342 19592 28122
rect 20372 27342 20382 28122
rect 19582 27332 19692 27342
rect 19682 26736 19692 27332
rect 19582 26726 19692 26736
rect 20272 27332 20382 27342
rect 20272 26736 20282 27332
rect 20272 26726 20382 26736
rect 19582 25946 19592 26726
rect 20372 25946 20382 26726
rect 19582 25936 19692 25946
rect 19160 25704 19408 25716
rect 19682 24784 19692 25936
rect 18876 24774 19692 24784
rect 20272 25936 20382 25946
rect 20272 24784 20282 25936
rect 20556 25716 20568 28256
rect 20792 25716 20804 28256
rect 21952 28256 22200 28718
rect 21078 28166 21678 28200
rect 21078 28132 21088 28166
rect 20978 28122 21088 28132
rect 21668 28132 21678 28166
rect 21668 28122 21778 28132
rect 20978 27342 20988 28122
rect 21768 27342 21778 28122
rect 20978 27332 21088 27342
rect 21078 26736 21088 27332
rect 20978 26726 21088 26736
rect 21668 27332 21778 27342
rect 21668 26736 21678 27332
rect 21668 26726 21778 26736
rect 20978 25946 20988 26726
rect 21768 25946 21778 26726
rect 20978 25936 21088 25946
rect 20556 25704 20804 25716
rect 21078 24784 21088 25936
rect 20272 24774 21088 24784
rect 21668 25936 21778 25946
rect 21668 24784 21678 25936
rect 21952 25716 21964 28256
rect 22188 25716 22200 28256
rect 23348 28256 23596 28718
rect 22474 28166 23074 28200
rect 22474 28132 22484 28166
rect 22374 28122 22484 28132
rect 23064 28132 23074 28166
rect 23064 28122 23174 28132
rect 22374 27342 22384 28122
rect 23164 27342 23174 28122
rect 22374 27332 22484 27342
rect 22474 26736 22484 27332
rect 22374 26726 22484 26736
rect 23064 27332 23174 27342
rect 23064 26736 23074 27332
rect 23064 26726 23174 26736
rect 22374 25946 22384 26726
rect 23164 25946 23174 26726
rect 22374 25936 22484 25946
rect 21952 25704 22200 25716
rect 22474 24784 22484 25936
rect 21668 24774 22484 24784
rect 23064 25936 23174 25946
rect 23064 24784 23074 25936
rect 23348 25716 23360 28256
rect 23584 25716 23596 28256
rect 24744 28256 24992 28718
rect 23870 28166 24470 28200
rect 23870 28132 23880 28166
rect 23770 28122 23880 28132
rect 24460 28132 24470 28166
rect 24460 28122 24570 28132
rect 23770 27342 23780 28122
rect 24560 27342 24570 28122
rect 23770 27332 23880 27342
rect 23870 26736 23880 27332
rect 23770 26726 23880 26736
rect 24460 27332 24570 27342
rect 24460 26736 24470 27332
rect 24460 26726 24570 26736
rect 23770 25946 23780 26726
rect 24560 25946 24570 26726
rect 23770 25936 23880 25946
rect 23348 25704 23596 25716
rect 23870 24784 23880 25936
rect 23064 24774 23880 24784
rect 24460 25936 24570 25946
rect 24460 24784 24470 25936
rect 24744 25716 24756 28256
rect 24980 25716 24992 28256
rect 26140 28256 26388 28718
rect 25266 28166 25866 28200
rect 25266 28132 25276 28166
rect 25166 28122 25276 28132
rect 25856 28132 25866 28166
rect 25856 28122 25966 28132
rect 25166 27342 25176 28122
rect 25956 27342 25966 28122
rect 25166 27332 25276 27342
rect 25266 26736 25276 27332
rect 25166 26726 25276 26736
rect 25856 27332 25966 27342
rect 25856 26736 25866 27332
rect 25856 26726 25966 26736
rect 25166 25946 25176 26726
rect 25956 25946 25966 26726
rect 25166 25936 25276 25946
rect 24744 25704 24992 25716
rect 25266 24784 25276 25936
rect 24460 24774 25276 24784
rect 25856 25936 25966 25946
rect 25856 24784 25866 25936
rect 26140 25716 26152 28256
rect 26376 25716 26388 28256
rect 27536 28256 27784 28718
rect 26662 28166 27262 28200
rect 26662 28132 26672 28166
rect 26562 28122 26672 28132
rect 27252 28132 27262 28166
rect 27252 28122 27362 28132
rect 26562 27342 26572 28122
rect 27352 27342 27362 28122
rect 26562 27332 26672 27342
rect 26662 26736 26672 27332
rect 26562 26726 26672 26736
rect 27252 27332 27362 27342
rect 27252 26736 27262 27332
rect 27252 26726 27362 26736
rect 26562 25946 26572 26726
rect 27352 25946 27362 26726
rect 26562 25936 26672 25946
rect 26140 25704 26388 25716
rect 26662 24784 26672 25936
rect 25856 24774 26672 24784
rect 27252 25936 27362 25946
rect 27252 24784 27262 25936
rect 27536 25716 27548 28256
rect 27772 25716 27784 28256
rect 28932 28256 29180 28718
rect 28058 28166 28658 28200
rect 28058 28132 28068 28166
rect 27958 28122 28068 28132
rect 28648 28132 28658 28166
rect 28648 28122 28758 28132
rect 27958 27342 27968 28122
rect 28748 27342 28758 28122
rect 27958 27332 28068 27342
rect 28058 26736 28068 27332
rect 27958 26726 28068 26736
rect 28648 27332 28758 27342
rect 28648 26736 28658 27332
rect 28648 26726 28758 26736
rect 27958 25946 27968 26726
rect 28748 25946 28758 26726
rect 27958 25936 28068 25946
rect 27536 25704 27784 25716
rect 28058 24784 28068 25936
rect 27252 24774 28068 24784
rect 28648 25936 28758 25946
rect 28648 24784 28658 25936
rect 28932 25716 28944 28256
rect 29168 25716 29180 28256
rect 30328 28256 30576 28718
rect 29454 28166 30054 28200
rect 29454 28132 29464 28166
rect 29352 28122 29464 28132
rect 30044 28132 30054 28166
rect 30044 28122 30154 28132
rect 29352 27342 29362 28122
rect 30144 27342 30154 28122
rect 29352 27332 29464 27342
rect 29454 26736 29464 27332
rect 29352 26726 29464 26736
rect 30044 27332 30154 27342
rect 30044 26736 30054 27332
rect 30044 26726 30154 26736
rect 29352 25946 29362 26726
rect 30144 25946 30154 26726
rect 29352 25936 29464 25946
rect 28932 25704 29180 25716
rect 29454 24784 29464 25936
rect 28648 24774 29464 24784
rect 30044 25936 30154 25946
rect 30044 24784 30054 25936
rect 30328 25716 30340 28256
rect 30564 25716 30576 28256
rect 31724 28256 31972 28718
rect 30850 28166 31450 28200
rect 30850 28132 30860 28166
rect 30750 28122 30860 28132
rect 31440 28132 31450 28166
rect 31440 28122 31550 28132
rect 30750 27342 30760 28122
rect 31540 27342 31550 28122
rect 30750 27332 30860 27342
rect 30850 26736 30860 27332
rect 30750 26726 30860 26736
rect 31440 27332 31550 27342
rect 31440 26736 31450 27332
rect 31440 26726 31550 26736
rect 30750 25946 30760 26726
rect 31540 25946 31550 26726
rect 30750 25936 30860 25946
rect 30328 25704 30576 25716
rect 30850 24784 30860 25936
rect 30044 24774 30860 24784
rect 31440 25936 31550 25946
rect 31440 24784 31450 25936
rect 31724 25716 31736 28256
rect 31960 25716 31972 28256
rect 33120 28256 33368 28718
rect 32246 28166 32846 28200
rect 32246 28132 32256 28166
rect 32146 28122 32256 28132
rect 32836 28132 32846 28166
rect 32836 28122 32946 28132
rect 32146 27342 32156 28122
rect 32936 27342 32946 28122
rect 32146 27332 32256 27342
rect 32246 26736 32256 27332
rect 32146 26726 32256 26736
rect 32836 27332 32946 27342
rect 32836 26736 32846 27332
rect 32836 26726 32946 26736
rect 32146 25946 32156 26726
rect 32936 25946 32946 26726
rect 32146 25936 32256 25946
rect 31724 25704 31972 25716
rect 32246 24784 32256 25936
rect 31440 24774 32256 24784
rect 32836 25936 32946 25946
rect 32836 24784 32846 25936
rect 33120 25716 33132 28256
rect 33356 25716 33368 28256
rect 34516 28256 34764 28718
rect 33642 28166 34242 28200
rect 33642 28132 33652 28166
rect 33542 28122 33652 28132
rect 34232 28132 34242 28166
rect 34232 28122 34342 28132
rect 33542 27342 33552 28122
rect 34332 27342 34342 28122
rect 33542 27332 33652 27342
rect 33642 26736 33652 27332
rect 33542 26726 33652 26736
rect 34232 27332 34342 27342
rect 34232 26736 34242 27332
rect 34232 26726 34342 26736
rect 33542 25946 33552 26726
rect 34332 25946 34342 26726
rect 33542 25936 33652 25946
rect 33120 25704 33368 25716
rect 33642 24784 33652 25936
rect 32836 24774 33652 24784
rect 34232 25936 34342 25946
rect 34232 24784 34242 25936
rect 34516 25716 34528 28256
rect 34752 25716 34764 28256
rect 35912 28256 36160 28718
rect 35038 28166 35638 28200
rect 35038 28132 35048 28166
rect 34938 28122 35048 28132
rect 35628 28132 35638 28166
rect 35628 28122 35738 28132
rect 34938 27342 34948 28122
rect 35728 27342 35738 28122
rect 34938 27332 35048 27342
rect 35038 26736 35048 27332
rect 34938 26726 35048 26736
rect 35628 27332 35738 27342
rect 35628 26736 35638 27332
rect 35628 26726 35738 26736
rect 34938 25946 34948 26726
rect 35728 25946 35738 26726
rect 34938 25936 35048 25946
rect 34516 25704 34764 25716
rect 35038 24784 35048 25936
rect 34232 24774 35048 24784
rect 35628 25936 35738 25946
rect 35628 24784 35638 25936
rect 35912 25716 35924 28256
rect 36148 25716 36160 28256
rect 37308 28256 37556 28718
rect 36434 28166 37034 28200
rect 36434 28132 36444 28166
rect 36334 28122 36444 28132
rect 37024 28132 37034 28166
rect 37024 28122 37134 28132
rect 36334 27342 36344 28122
rect 37124 27342 37134 28122
rect 36334 27332 36444 27342
rect 36434 26736 36444 27332
rect 36334 26726 36444 26736
rect 37024 27332 37134 27342
rect 37024 26736 37034 27332
rect 37024 26726 37134 26736
rect 36334 25946 36344 26726
rect 37124 25946 37134 26726
rect 36334 25936 36444 25946
rect 35912 25704 36160 25716
rect 36434 24784 36444 25936
rect 35628 24774 36444 24784
rect 37024 25936 37134 25946
rect 37024 24784 37034 25936
rect 37308 25716 37320 28256
rect 37544 25716 37556 28256
rect 38704 28256 38952 28718
rect 37830 28166 38430 28200
rect 37830 28132 37840 28166
rect 37730 28122 37840 28132
rect 38420 28132 38430 28166
rect 38420 28122 38530 28132
rect 37730 27342 37740 28122
rect 38520 27342 38530 28122
rect 37730 27332 37840 27342
rect 37830 26736 37840 27332
rect 37730 26726 37840 26736
rect 38420 27332 38530 27342
rect 38420 26736 38430 27332
rect 38420 26726 38530 26736
rect 37730 25946 37740 26726
rect 38520 25946 38530 26726
rect 37730 25936 37840 25946
rect 37308 25704 37556 25716
rect 37830 24784 37840 25936
rect 37024 24774 37840 24784
rect 38420 25936 38530 25946
rect 38420 24784 38430 25936
rect 38704 25716 38716 28256
rect 38940 25716 38952 28256
rect 40100 28256 40348 28718
rect 39226 28166 39826 28200
rect 39226 28132 39236 28166
rect 39126 28122 39236 28132
rect 39816 28132 39826 28166
rect 39816 28122 39926 28132
rect 39126 27342 39136 28122
rect 39916 27342 39926 28122
rect 39126 27332 39236 27342
rect 39226 26736 39236 27332
rect 39126 26726 39236 26736
rect 39816 27332 39926 27342
rect 39816 26736 39826 27332
rect 39816 26726 39926 26736
rect 39126 25946 39136 26726
rect 39916 25946 39926 26726
rect 39126 25936 39236 25946
rect 38704 25704 38952 25716
rect 39226 24784 39236 25936
rect 38420 24774 39236 24784
rect 39816 25936 39926 25946
rect 39816 24784 39826 25936
rect 40100 25716 40112 28256
rect 40336 25716 40348 28256
rect 41496 28256 41744 28718
rect 40622 28166 41222 28200
rect 40622 28132 40632 28166
rect 40522 28122 40632 28132
rect 41212 28132 41222 28166
rect 41212 28122 41322 28132
rect 40522 27342 40532 28122
rect 41312 27342 41322 28122
rect 40522 27332 40632 27342
rect 40622 26736 40632 27332
rect 40522 26726 40632 26736
rect 41212 27332 41322 27342
rect 41212 26736 41222 27332
rect 41212 26726 41322 26736
rect 40522 25946 40532 26726
rect 41312 25946 41322 26726
rect 40522 25936 40632 25946
rect 40100 25704 40348 25716
rect 40622 24784 40632 25936
rect 39816 24774 40632 24784
rect 41212 25936 41322 25946
rect 41212 24784 41222 25936
rect 41496 25716 41508 28256
rect 41732 25716 41744 28256
rect 42892 28256 43140 28718
rect 42018 28166 42618 28200
rect 42018 28132 42028 28166
rect 41918 28122 42028 28132
rect 42608 28132 42618 28166
rect 42608 28122 42718 28132
rect 41918 27342 41928 28122
rect 42708 27342 42718 28122
rect 41918 27332 42028 27342
rect 42018 26736 42028 27332
rect 41918 26726 42028 26736
rect 42608 27332 42718 27342
rect 42608 26736 42618 27332
rect 42608 26726 42718 26736
rect 41918 25946 41928 26726
rect 42708 25946 42718 26726
rect 41918 25936 42028 25946
rect 41496 25704 41744 25716
rect 42018 24784 42028 25936
rect 41212 24774 42028 24784
rect 42608 25936 42718 25946
rect 42608 24784 42618 25936
rect 42892 25716 42904 28256
rect 43128 25716 43140 28256
rect 44288 28256 44536 28718
rect 43414 28166 44014 28200
rect 43414 28132 43424 28166
rect 43314 28122 43424 28132
rect 44004 28132 44014 28166
rect 44004 28122 44114 28132
rect 43314 27342 43324 28122
rect 44104 27342 44114 28122
rect 43314 27332 43424 27342
rect 43414 26736 43424 27332
rect 43314 26726 43424 26736
rect 44004 27332 44114 27342
rect 44004 26736 44014 27332
rect 44004 26726 44114 26736
rect 43314 25946 43324 26726
rect 44104 25946 44114 26726
rect 43314 25936 43424 25946
rect 42892 25704 43140 25716
rect 43414 24784 43424 25936
rect 42608 24774 43424 24784
rect 44004 25936 44114 25946
rect 44004 24784 44014 25936
rect 44288 25716 44300 28256
rect 44524 25716 44536 28256
rect 45684 28256 45932 28718
rect 44810 28166 45410 28200
rect 44810 28132 44820 28166
rect 44710 28122 44820 28132
rect 45400 28132 45410 28166
rect 45400 28122 45510 28132
rect 44710 27342 44720 28122
rect 45500 27342 45510 28122
rect 44710 27332 44820 27342
rect 44810 26736 44820 27332
rect 44710 26726 44820 26736
rect 45400 27332 45510 27342
rect 45400 26736 45410 27332
rect 45400 26726 45510 26736
rect 44710 25946 44720 26726
rect 45500 25946 45510 26726
rect 44710 25936 44820 25946
rect 44288 25704 44536 25716
rect 44810 24784 44820 25936
rect 44004 24774 44820 24784
rect 45400 25936 45510 25946
rect 45400 24784 45410 25936
rect 45684 25716 45696 28256
rect 45920 25716 45932 28256
rect 47080 28256 47328 28718
rect 46206 28166 46806 28200
rect 46206 28132 46216 28166
rect 46106 28122 46216 28132
rect 46796 28132 46806 28166
rect 46796 28122 46906 28132
rect 46106 27342 46116 28122
rect 46896 27342 46906 28122
rect 46106 27332 46216 27342
rect 46206 26736 46216 27332
rect 46106 26726 46216 26736
rect 46796 27332 46906 27342
rect 46796 26736 46806 27332
rect 46796 26726 46906 26736
rect 46106 25946 46116 26726
rect 46896 25946 46906 26726
rect 46106 25936 46216 25946
rect 45684 25704 45932 25716
rect 46206 24784 46216 25936
rect 45400 24774 46216 24784
rect 46796 25936 46906 25946
rect 46796 24784 46806 25936
rect 47080 25716 47092 28256
rect 47316 25716 47328 28256
rect 48476 28256 48724 28718
rect 47602 28166 48202 28200
rect 47602 28132 47612 28166
rect 47502 28122 47612 28132
rect 48192 28132 48202 28166
rect 48192 28122 48302 28132
rect 47502 27342 47512 28122
rect 48292 27342 48302 28122
rect 47502 27332 47612 27342
rect 47602 26736 47612 27332
rect 47502 26726 47612 26736
rect 48192 27332 48302 27342
rect 48192 26736 48202 27332
rect 48192 26726 48302 26736
rect 47502 25946 47512 26726
rect 48292 25946 48302 26726
rect 47502 25936 47612 25946
rect 47080 25704 47328 25716
rect 47602 24784 47612 25936
rect 46796 24774 47612 24784
rect 48192 25936 48302 25946
rect 48192 24784 48202 25936
rect 48476 25716 48488 28256
rect 48712 25716 48724 28256
rect 49872 28256 50120 28718
rect 48998 28166 49598 28200
rect 48998 28132 49008 28166
rect 48898 28122 49008 28132
rect 49588 28132 49598 28166
rect 49588 28122 49698 28132
rect 48898 27342 48908 28122
rect 49688 27342 49698 28122
rect 48898 27332 49008 27342
rect 48998 26736 49008 27332
rect 48898 26726 49008 26736
rect 49588 27332 49698 27342
rect 49588 26736 49598 27332
rect 49588 26726 49698 26736
rect 48898 25946 48908 26726
rect 49688 25946 49698 26726
rect 48898 25936 49008 25946
rect 48476 25704 48724 25716
rect 48998 24784 49008 25936
rect 48192 24774 49008 24784
rect 49588 25936 49698 25946
rect 49588 24784 49598 25936
rect 49872 25716 49884 28256
rect 50108 25716 50120 28256
rect 50394 28166 50994 28200
rect 50394 28132 50404 28166
rect 50294 28122 50404 28132
rect 50984 28132 50994 28166
rect 50984 28122 51094 28132
rect 50294 27342 50304 28122
rect 51084 27342 51094 28122
rect 50294 27332 50404 27342
rect 50394 26736 50404 27332
rect 50294 26726 50404 26736
rect 50984 27332 51094 27342
rect 50984 26736 50994 27332
rect 50984 26726 51094 26736
rect 50294 25946 50304 26726
rect 51084 25946 51094 26726
rect 50294 25936 50404 25946
rect 49872 25704 50120 25716
rect 50394 24784 50404 25936
rect 49588 24774 50404 24784
rect 50984 25936 51094 25946
rect 50984 24784 50994 25936
rect 50984 24774 70094 24784
rect -2992 24438 3654 24448
rect -2992 23856 -1228 24438
rect 3618 23856 3654 24438
rect 4632 24394 4642 24774
rect 70084 24394 70094 24774
rect 4632 24384 70094 24394
rect 4632 24284 4680 24384
rect 4948 24284 4996 24384
rect 5264 24284 5312 24384
rect 5580 24284 5628 24384
rect 5896 24284 5944 24384
rect 6212 24284 6260 24384
rect 6528 24284 6576 24384
rect 6844 24284 6892 24384
rect 7160 24284 7208 24384
rect 7476 24284 7524 24384
rect 7792 24284 7840 24384
rect 8108 24284 8156 24384
rect 8424 24284 8472 24384
rect 8740 24284 8788 24384
rect 9056 24284 9104 24384
rect 9372 24284 9420 24384
rect 9688 24284 9736 24384
rect 10004 24284 10052 24384
rect 10320 24284 10368 24384
rect 10636 24284 10684 24384
rect 10952 24284 11000 24384
rect 11268 24284 11316 24384
rect 11584 24284 11632 24384
rect 11900 24284 11948 24384
rect 12216 24284 12264 24384
rect 12532 24284 12580 24384
rect 12848 24284 12896 24384
rect 13164 24284 13212 24384
rect 13480 24284 13528 24384
rect 13796 24284 13844 24384
rect 14112 24284 14160 24384
rect 14428 24284 14476 24384
rect 14744 24284 14792 24384
rect 15060 24284 15108 24384
rect 15376 24284 15424 24384
rect 15692 24284 15740 24384
rect 16008 24284 16056 24384
rect 16324 24284 16372 24384
rect 16640 24284 16688 24384
rect 16956 24284 17004 24384
rect 17272 24284 17320 24384
rect 17786 24284 17834 24384
rect 18102 24284 18150 24384
rect 18418 24284 18466 24384
rect 18734 24284 18782 24384
rect 19050 24284 19098 24384
rect 19366 24284 19414 24384
rect 19682 24284 19730 24384
rect 19998 24284 20046 24384
rect 20314 24284 20362 24384
rect 20630 24284 20678 24384
rect 20946 24284 20994 24384
rect 21262 24284 21310 24384
rect 21578 24284 21626 24384
rect 21894 24284 21942 24384
rect 22210 24284 22258 24384
rect 22526 24284 22574 24384
rect 22842 24284 22890 24384
rect 23158 24284 23206 24384
rect 23474 24284 23522 24384
rect 23790 24284 23838 24384
rect 24106 24284 24154 24384
rect 24422 24284 24470 24384
rect 24738 24284 24786 24384
rect 25054 24284 25102 24384
rect 25370 24284 25418 24384
rect 25686 24284 25734 24384
rect 26002 24284 26050 24384
rect 26318 24284 26366 24384
rect 26634 24284 26682 24384
rect 26950 24284 26998 24384
rect 27266 24284 27314 24384
rect 27582 24284 27630 24384
rect 27898 24284 27946 24384
rect 28214 24284 28262 24384
rect 28530 24284 28578 24384
rect 28846 24284 28894 24384
rect 29162 24284 29210 24384
rect 29478 24284 29526 24384
rect 29794 24284 29842 24384
rect 30110 24284 30158 24384
rect 30426 24284 30474 24384
rect 30940 24284 30988 24384
rect 31256 24284 31304 24384
rect 31572 24284 31620 24384
rect 31888 24284 31936 24384
rect 32204 24284 32252 24384
rect 32520 24284 32568 24384
rect 32836 24284 32884 24384
rect 33152 24284 33200 24384
rect 33468 24284 33516 24384
rect 33784 24284 33832 24384
rect 34100 24284 34148 24384
rect 34416 24284 34464 24384
rect 34732 24284 34780 24384
rect 35048 24284 35096 24384
rect 35364 24284 35412 24384
rect 35680 24284 35728 24384
rect 35996 24284 36044 24384
rect 36312 24284 36360 24384
rect 36628 24284 36676 24384
rect 36944 24284 36992 24384
rect 37260 24284 37308 24384
rect 37576 24284 37624 24384
rect 37892 24284 37940 24384
rect 38208 24284 38256 24384
rect 38524 24284 38572 24384
rect 38840 24284 38888 24384
rect 39156 24284 39204 24384
rect 39472 24284 39520 24384
rect 39788 24284 39836 24384
rect 40104 24284 40152 24384
rect 40420 24284 40468 24384
rect 40736 24284 40784 24384
rect 41052 24284 41100 24384
rect 41368 24284 41416 24384
rect 41684 24284 41732 24384
rect 42000 24284 42048 24384
rect 42316 24284 42364 24384
rect 42632 24284 42680 24384
rect 42948 24284 42996 24384
rect 43264 24284 43312 24384
rect 43580 24284 43628 24384
rect 44094 24284 44142 24384
rect 44410 24284 44458 24384
rect 44726 24284 44774 24384
rect 45042 24284 45090 24384
rect 45358 24284 45406 24384
rect 45674 24284 45722 24384
rect 45990 24284 46038 24384
rect 46306 24284 46354 24384
rect 46622 24284 46670 24384
rect 46938 24284 46986 24384
rect 47254 24284 47302 24384
rect 47570 24284 47618 24384
rect 47886 24284 47934 24384
rect 48202 24284 48250 24384
rect 48518 24284 48566 24384
rect 48834 24284 48882 24384
rect 49150 24284 49198 24384
rect 49466 24284 49514 24384
rect 49782 24284 49830 24384
rect 50098 24284 50146 24384
rect 50414 24284 50462 24384
rect 50730 24284 50778 24384
rect 51046 24284 51094 24384
rect 51362 24284 51410 24384
rect 51678 24284 51726 24384
rect 51994 24284 52042 24384
rect 52310 24284 52358 24384
rect 52626 24284 52674 24384
rect 52942 24284 52990 24384
rect 53258 24284 53306 24384
rect 53574 24284 53622 24384
rect 53890 24284 53938 24384
rect 54206 24284 54254 24384
rect 54522 24284 54570 24384
rect 54838 24284 54886 24384
rect 55154 24284 55202 24384
rect 55470 24284 55518 24384
rect 55786 24284 55834 24384
rect 56102 24284 56150 24384
rect 56418 24284 56466 24384
rect 56734 24284 56782 24384
rect 57248 24284 57296 24384
rect 57564 24284 57612 24384
rect 57880 24284 57928 24384
rect 58196 24284 58244 24384
rect 58512 24284 58560 24384
rect 58828 24284 58876 24384
rect 59144 24284 59192 24384
rect 59460 24284 59508 24384
rect 59776 24284 59824 24384
rect 60092 24284 60140 24384
rect 60408 24284 60456 24384
rect 60724 24284 60772 24384
rect 61040 24284 61088 24384
rect 61356 24284 61404 24384
rect 61672 24284 61720 24384
rect 61988 24284 62036 24384
rect 62304 24284 62352 24384
rect 62620 24284 62668 24384
rect 62936 24284 62984 24384
rect 63252 24284 63300 24384
rect 63568 24284 63616 24384
rect 63884 24284 63932 24384
rect 64200 24284 64248 24384
rect 64516 24284 64564 24384
rect 64832 24284 64880 24384
rect 65148 24284 65196 24384
rect 65464 24284 65512 24384
rect 65780 24284 65828 24384
rect 66096 24284 66144 24384
rect 66412 24284 66460 24384
rect 66728 24284 66776 24384
rect 67044 24284 67092 24384
rect 67360 24284 67408 24384
rect 67676 24284 67724 24384
rect 67992 24284 68040 24384
rect 68308 24284 68356 24384
rect 68624 24284 68672 24384
rect 68940 24284 68988 24384
rect 69256 24284 69304 24384
rect 69572 24284 69620 24384
rect 69888 24284 69936 24384
rect -2992 23846 3654 23856
rect 3690 23336 4106 23344
rect 3690 22936 3698 23336
rect 4098 22936 4106 23336
rect 3690 22928 4106 22936
rect -2980 19040 -2560 19048
rect -2980 18640 -2968 19040
rect -2568 18640 -2560 19040
rect -2980 18630 -2560 18640
rect 4790 14276 4838 14372
rect 5106 14276 5154 14372
rect 5422 14276 5470 14372
rect 5738 14276 5786 14372
rect 6054 14276 6102 14372
rect 6370 14276 6418 14372
rect 6686 14276 6734 14372
rect 7002 14276 7050 14372
rect 7318 14276 7366 14372
rect 7634 14276 7682 14372
rect 7950 14276 7998 14372
rect 8266 14276 8314 14372
rect 8582 14276 8630 14372
rect 8898 14276 8946 14372
rect 9214 14276 9262 14372
rect 9530 14276 9578 14372
rect 9846 14276 9894 14372
rect 10162 14276 10210 14372
rect 10478 14276 10526 14372
rect 10794 14276 10842 14372
rect 11110 14276 11158 14372
rect 11426 14276 11474 14372
rect 11742 14276 11790 14372
rect 12058 14276 12106 14372
rect 12374 14276 12422 14372
rect 12690 14276 12738 14372
rect 13006 14276 13054 14372
rect 13322 14276 13370 14372
rect 13638 14276 13686 14372
rect 13954 14276 14002 14372
rect 14270 14276 14318 14372
rect 14586 14276 14634 14372
rect 14902 14276 14950 14372
rect 15218 14276 15266 14372
rect 15534 14276 15582 14372
rect 15850 14276 15898 14372
rect 16166 14276 16214 14372
rect 16482 14276 16530 14372
rect 16798 14276 16846 14372
rect 17114 14276 17162 14372
rect 17944 14276 17992 14372
rect 18260 14276 18308 14372
rect 18576 14276 18624 14372
rect 18892 14276 18940 14372
rect 19208 14276 19256 14372
rect 19524 14276 19572 14372
rect 19840 14276 19888 14372
rect 20156 14276 20204 14372
rect 20472 14276 20520 14372
rect 20788 14276 20836 14372
rect 21104 14276 21152 14372
rect 21420 14276 21468 14372
rect 21736 14276 21784 14372
rect 22052 14276 22100 14372
rect 22368 14276 22416 14372
rect 22684 14276 22732 14372
rect 23000 14276 23048 14372
rect 23316 14276 23364 14372
rect 23632 14276 23680 14372
rect 23948 14276 23996 14372
rect 24264 14276 24312 14372
rect 24580 14276 24628 14372
rect 24896 14276 24944 14372
rect 25212 14276 25260 14372
rect 25528 14276 25576 14372
rect 25844 14276 25892 14372
rect 26160 14276 26208 14372
rect 26476 14276 26524 14372
rect 26792 14276 26840 14372
rect 27108 14276 27156 14372
rect 27424 14276 27472 14372
rect 27740 14276 27788 14372
rect 28056 14276 28104 14372
rect 28372 14276 28420 14372
rect 28688 14276 28736 14372
rect 29004 14276 29052 14372
rect 29320 14276 29368 14372
rect 29636 14276 29684 14372
rect 29952 14276 30000 14372
rect 30268 14276 30316 14372
rect 31098 14276 31146 14372
rect 31414 14276 31462 14372
rect 31730 14276 31778 14372
rect 32046 14276 32094 14372
rect 32362 14276 32410 14372
rect 32678 14276 32726 14372
rect 32994 14276 33042 14372
rect 33310 14276 33358 14372
rect 33626 14276 33674 14372
rect 33942 14276 33990 14372
rect 34258 14276 34306 14372
rect 34574 14276 34622 14372
rect 34890 14276 34938 14372
rect 35206 14276 35254 14372
rect 35522 14276 35570 14372
rect 35838 14276 35886 14372
rect 36154 14276 36202 14372
rect 36470 14276 36518 14372
rect 36786 14276 36834 14372
rect 37102 14276 37150 14372
rect 37418 14276 37466 14372
rect 37734 14276 37782 14372
rect 38050 14276 38098 14372
rect 38366 14276 38414 14372
rect 38682 14276 38730 14372
rect 38998 14276 39046 14372
rect 39314 14276 39362 14372
rect 39630 14276 39678 14372
rect 39946 14276 39994 14372
rect 40262 14276 40310 14372
rect 40578 14276 40626 14372
rect 40894 14276 40942 14372
rect 41210 14276 41258 14372
rect 41526 14276 41574 14372
rect 41842 14276 41890 14372
rect 42158 14276 42206 14372
rect 42474 14276 42522 14372
rect 42790 14276 42838 14372
rect 43106 14276 43154 14372
rect 43422 14276 43470 14372
rect 44252 14276 44300 14372
rect 44568 14276 44616 14372
rect 44884 14276 44932 14372
rect 45200 14276 45248 14372
rect 45516 14276 45564 14372
rect 45832 14276 45880 14372
rect 46148 14276 46196 14372
rect 46464 14276 46512 14372
rect 46780 14276 46828 14372
rect 47096 14276 47144 14372
rect 47412 14276 47460 14372
rect 47728 14276 47776 14372
rect 48044 14276 48092 14372
rect 48360 14276 48408 14372
rect 48676 14276 48724 14372
rect 48992 14276 49040 14372
rect 49308 14276 49356 14372
rect 49624 14276 49672 14372
rect 49940 14276 49988 14372
rect 50256 14276 50304 14372
rect 50572 14276 50620 14372
rect 50888 14276 50936 14372
rect 51204 14276 51252 14372
rect 51520 14276 51568 14372
rect 51836 14276 51884 14372
rect 52152 14276 52200 14372
rect 52468 14276 52516 14372
rect 52784 14276 52832 14372
rect 53100 14276 53148 14372
rect 53416 14276 53464 14372
rect 53732 14276 53780 14372
rect 54048 14276 54096 14372
rect 54364 14276 54412 14372
rect 54680 14276 54728 14372
rect 54996 14276 55044 14372
rect 55312 14276 55360 14372
rect 55628 14276 55676 14372
rect 55944 14276 55992 14372
rect 56260 14276 56308 14372
rect 56576 14276 56624 14372
rect 57406 14276 57454 14372
rect 57722 14276 57770 14372
rect 58038 14276 58086 14372
rect 58354 14276 58402 14372
rect 58670 14276 58718 14372
rect 58986 14276 59034 14372
rect 59302 14276 59350 14372
rect 59618 14276 59666 14372
rect 59934 14276 59982 14372
rect 60250 14276 60298 14372
rect 60566 14276 60614 14372
rect 60882 14276 60930 14372
rect 61198 14276 61246 14372
rect 61514 14276 61562 14372
rect 61830 14276 61878 14372
rect 62146 14276 62194 14372
rect 62462 14276 62510 14372
rect 62778 14276 62826 14372
rect 63094 14276 63142 14372
rect 63410 14276 63458 14372
rect 63726 14276 63774 14372
rect 64042 14276 64090 14372
rect 64358 14276 64406 14372
rect 64674 14276 64722 14372
rect 64990 14276 65038 14372
rect 65306 14276 65354 14372
rect 65622 14276 65670 14372
rect 65938 14276 65986 14372
rect 66254 14276 66302 14372
rect 66570 14276 66618 14372
rect 66886 14276 66934 14372
rect 67202 14276 67250 14372
rect 67518 14276 67566 14372
rect 67834 14276 67882 14372
rect 68150 14276 68198 14372
rect 68466 14276 68514 14372
rect 68782 14276 68830 14372
rect 69098 14276 69146 14372
rect 69414 14276 69462 14372
rect 69730 14276 69778 14372
rect 4568 14182 69954 14276
rect 526 13434 3458 13438
rect 526 13426 3460 13434
rect 526 13370 538 13426
rect 3448 13370 3460 13426
rect 526 13360 3460 13370
rect 526 13358 616 13360
rect 842 13358 932 13360
rect 1158 13358 1248 13360
rect 1474 13358 1564 13360
rect 1790 13358 1880 13360
rect 2106 13358 2196 13360
rect 2422 13358 2512 13360
rect 2738 13358 2828 13360
rect 3054 13358 3144 13360
rect 3370 13358 3460 13360
rect -13830 4844 -13230 12596
rect -11792 11568 -5364 11888
rect -12170 11332 -11950 11356
rect -12170 10956 -12146 11332
rect -11974 10956 -11950 11332
rect -12170 9726 -11950 10956
rect -12170 9350 -12146 9726
rect -11974 9350 -11950 9726
rect -12170 8120 -11950 9350
rect -12170 7744 -12146 8120
rect -11974 7744 -11950 8120
rect -12170 6514 -11950 7744
rect -12170 6138 -12146 6514
rect -11974 6138 -11950 6514
rect -12170 5264 -11950 6138
rect -11792 10854 -11786 11568
rect -11586 11528 -10380 11568
rect -11586 10854 -11580 11528
rect -11792 9962 -11580 10854
rect -11792 9114 -11786 9962
rect -11586 9114 -11580 9962
rect -11792 8356 -11580 9114
rect -11792 7508 -11786 8356
rect -11586 7508 -11580 8356
rect -11792 6750 -11580 7508
rect -11792 5902 -11786 6750
rect -11586 5902 -11580 6750
rect -11792 5884 -11580 5902
rect -10764 11332 -10544 11356
rect -10764 10956 -10740 11332
rect -10568 10956 -10544 11332
rect -10764 9726 -10544 10956
rect -10764 9350 -10740 9726
rect -10568 9350 -10544 9726
rect -10764 8120 -10544 9350
rect -10764 7744 -10740 8120
rect -10568 7744 -10544 8120
rect -10764 6514 -10544 7744
rect -10764 6138 -10740 6514
rect -10568 6138 -10544 6514
rect -10764 5264 -10544 6138
rect -10386 10854 -10380 11528
rect -10180 11528 -8974 11568
rect -10180 10854 -10174 11528
rect -10386 9962 -10174 10854
rect -10386 9114 -10380 9962
rect -10180 9114 -10174 9962
rect -10386 8356 -10174 9114
rect -10386 7508 -10380 8356
rect -10180 7508 -10174 8356
rect -10386 6750 -10174 7508
rect -10386 5902 -10380 6750
rect -10180 5902 -10174 6750
rect -10386 5884 -10174 5902
rect -9358 11332 -9138 11356
rect -9358 10956 -9334 11332
rect -9162 10956 -9138 11332
rect -9358 9726 -9138 10956
rect -9358 9350 -9334 9726
rect -9162 9350 -9138 9726
rect -9358 8120 -9138 9350
rect -9358 7744 -9334 8120
rect -9162 7744 -9138 8120
rect -9358 6514 -9138 7744
rect -9358 6138 -9334 6514
rect -9162 6138 -9138 6514
rect -9358 5264 -9138 6138
rect -8980 10854 -8974 11528
rect -8774 11528 -7568 11568
rect -8774 10854 -8768 11528
rect -8980 9962 -8768 10854
rect -8980 9114 -8974 9962
rect -8774 9114 -8768 9962
rect -8980 8356 -8768 9114
rect -8980 7508 -8974 8356
rect -8774 7508 -8768 8356
rect -8980 6750 -8768 7508
rect -8980 5902 -8974 6750
rect -8774 5902 -8768 6750
rect -8980 5884 -8768 5902
rect -7952 11332 -7732 11356
rect -7952 10956 -7928 11332
rect -7756 10956 -7732 11332
rect -7952 9726 -7732 10956
rect -7952 9350 -7928 9726
rect -7756 9350 -7732 9726
rect -7952 8120 -7732 9350
rect -7952 7744 -7928 8120
rect -7756 7744 -7732 8120
rect -7952 6514 -7732 7744
rect -7952 6138 -7928 6514
rect -7756 6138 -7732 6514
rect -7952 5264 -7732 6138
rect -7574 10854 -7568 11528
rect -7368 11528 -5364 11568
rect -7368 10854 -7362 11528
rect -7574 9962 -7362 10854
rect -7574 9114 -7568 9962
rect -7368 9114 -7362 9962
rect -7574 8356 -7362 9114
rect -5724 9254 -5364 11528
rect -3880 11686 -3870 12886
rect -3290 11686 -3280 12886
rect -3880 11676 -3280 11686
rect -3880 11088 -3280 11094
rect 540 13202 606 13358
rect 540 13004 546 13202
rect 600 13004 606 13202
rect 540 12890 606 13004
rect 540 12692 546 12890
rect 600 12692 606 12890
rect 540 12578 606 12692
rect 540 12386 546 12578
rect 600 12386 606 12578
rect 540 12268 606 12386
rect 540 12076 546 12268
rect 598 12076 606 12268
rect 540 11958 606 12076
rect 540 11766 546 11958
rect 598 11766 606 11958
rect 540 11644 606 11766
rect 540 11456 546 11644
rect 598 11456 606 11644
rect 540 11334 606 11456
rect 540 11146 546 11334
rect 598 11146 606 11334
rect 540 11026 606 11146
rect 540 10838 546 11026
rect 598 10838 606 11026
rect 540 10712 606 10838
rect 540 10526 546 10712
rect 598 10526 606 10712
rect 540 10404 606 10526
rect 540 10218 546 10404
rect 598 10218 606 10404
rect 540 10060 606 10218
rect 856 13202 922 13358
rect 856 13004 862 13202
rect 916 13004 922 13202
rect 856 12890 922 13004
rect 856 12692 862 12890
rect 916 12692 922 12890
rect 856 12578 922 12692
rect 856 12386 862 12578
rect 916 12386 922 12578
rect 856 12268 922 12386
rect 856 12076 862 12268
rect 914 12076 922 12268
rect 856 11958 922 12076
rect 856 11766 862 11958
rect 914 11766 922 11958
rect 856 11644 922 11766
rect 856 11456 862 11644
rect 914 11456 922 11644
rect 856 11334 922 11456
rect 856 11146 862 11334
rect 914 11146 922 11334
rect 856 11026 922 11146
rect 856 10838 862 11026
rect 914 10838 922 11026
rect 856 10712 922 10838
rect 856 10526 862 10712
rect 914 10526 922 10712
rect 856 10404 922 10526
rect 856 10218 862 10404
rect 914 10218 922 10404
rect 856 10060 922 10218
rect 1172 13202 1238 13358
rect 1172 13004 1178 13202
rect 1232 13004 1238 13202
rect 1172 12890 1238 13004
rect 1172 12692 1178 12890
rect 1232 12692 1238 12890
rect 1172 12578 1238 12692
rect 1172 12386 1178 12578
rect 1232 12386 1238 12578
rect 1172 12268 1238 12386
rect 1172 12076 1178 12268
rect 1230 12076 1238 12268
rect 1172 11958 1238 12076
rect 1172 11766 1178 11958
rect 1230 11766 1238 11958
rect 1172 11644 1238 11766
rect 1172 11456 1178 11644
rect 1230 11456 1238 11644
rect 1172 11334 1238 11456
rect 1172 11146 1178 11334
rect 1230 11146 1238 11334
rect 1172 11026 1238 11146
rect 1172 10838 1178 11026
rect 1230 10838 1238 11026
rect 1172 10712 1238 10838
rect 1172 10526 1178 10712
rect 1230 10526 1238 10712
rect 1172 10404 1238 10526
rect 1172 10218 1178 10404
rect 1230 10218 1238 10404
rect 1172 10060 1238 10218
rect 1488 13202 1554 13358
rect 1488 13004 1494 13202
rect 1548 13004 1554 13202
rect 1488 12890 1554 13004
rect 1488 12692 1494 12890
rect 1548 12692 1554 12890
rect 1488 12578 1554 12692
rect 1488 12386 1494 12578
rect 1548 12386 1554 12578
rect 1488 12268 1554 12386
rect 1488 12076 1494 12268
rect 1546 12076 1554 12268
rect 1488 11958 1554 12076
rect 1488 11766 1494 11958
rect 1546 11766 1554 11958
rect 1488 11644 1554 11766
rect 1488 11456 1494 11644
rect 1546 11456 1554 11644
rect 1488 11334 1554 11456
rect 1488 11146 1494 11334
rect 1546 11146 1554 11334
rect 1488 11026 1554 11146
rect 1488 10838 1494 11026
rect 1546 10838 1554 11026
rect 1488 10712 1554 10838
rect 1488 10526 1494 10712
rect 1546 10526 1554 10712
rect 1488 10404 1554 10526
rect 1488 10218 1494 10404
rect 1546 10218 1554 10404
rect 1488 10060 1554 10218
rect 1804 13202 1870 13358
rect 1804 13004 1810 13202
rect 1864 13004 1870 13202
rect 1804 12890 1870 13004
rect 1804 12692 1810 12890
rect 1864 12692 1870 12890
rect 1804 12578 1870 12692
rect 1804 12386 1810 12578
rect 1864 12386 1870 12578
rect 1804 12268 1870 12386
rect 1804 12076 1810 12268
rect 1862 12076 1870 12268
rect 1804 11958 1870 12076
rect 1804 11766 1810 11958
rect 1862 11766 1870 11958
rect 1804 11644 1870 11766
rect 1804 11456 1810 11644
rect 1862 11456 1870 11644
rect 1804 11334 1870 11456
rect 1804 11146 1810 11334
rect 1862 11146 1870 11334
rect 1804 11026 1870 11146
rect 1804 10838 1810 11026
rect 1862 10838 1870 11026
rect 1804 10712 1870 10838
rect 1804 10526 1810 10712
rect 1862 10526 1870 10712
rect 1804 10404 1870 10526
rect 1804 10218 1810 10404
rect 1862 10218 1870 10404
rect 1804 10060 1870 10218
rect 2120 13202 2186 13358
rect 2120 13004 2126 13202
rect 2180 13004 2186 13202
rect 2120 12890 2186 13004
rect 2120 12692 2126 12890
rect 2180 12692 2186 12890
rect 2120 12578 2186 12692
rect 2120 12386 2126 12578
rect 2180 12386 2186 12578
rect 2120 12268 2186 12386
rect 2120 12076 2126 12268
rect 2178 12076 2186 12268
rect 2120 11958 2186 12076
rect 2120 11766 2126 11958
rect 2178 11766 2186 11958
rect 2120 11644 2186 11766
rect 2120 11456 2126 11644
rect 2178 11456 2186 11644
rect 2120 11334 2186 11456
rect 2120 11146 2126 11334
rect 2178 11146 2186 11334
rect 2120 11026 2186 11146
rect 2120 10838 2126 11026
rect 2178 10838 2186 11026
rect 2120 10712 2186 10838
rect 2120 10526 2126 10712
rect 2178 10526 2186 10712
rect 2120 10404 2186 10526
rect 2120 10218 2126 10404
rect 2178 10218 2186 10404
rect 2120 10060 2186 10218
rect 2436 13202 2502 13358
rect 2436 13004 2442 13202
rect 2496 13004 2502 13202
rect 2436 12890 2502 13004
rect 2436 12692 2442 12890
rect 2496 12692 2502 12890
rect 2436 12578 2502 12692
rect 2436 12386 2442 12578
rect 2496 12386 2502 12578
rect 2436 12268 2502 12386
rect 2436 12076 2442 12268
rect 2494 12076 2502 12268
rect 2436 11958 2502 12076
rect 2436 11766 2442 11958
rect 2494 11766 2502 11958
rect 2436 11644 2502 11766
rect 2436 11456 2442 11644
rect 2494 11456 2502 11644
rect 2436 11334 2502 11456
rect 2436 11146 2442 11334
rect 2494 11146 2502 11334
rect 2436 11026 2502 11146
rect 2436 10838 2442 11026
rect 2494 10838 2502 11026
rect 2436 10712 2502 10838
rect 2436 10526 2442 10712
rect 2494 10526 2502 10712
rect 2436 10404 2502 10526
rect 2436 10218 2442 10404
rect 2494 10218 2502 10404
rect 2436 10060 2502 10218
rect 2752 13202 2818 13358
rect 2752 13004 2758 13202
rect 2812 13004 2818 13202
rect 2752 12890 2818 13004
rect 2752 12692 2758 12890
rect 2812 12692 2818 12890
rect 2752 12578 2818 12692
rect 2752 12386 2758 12578
rect 2812 12386 2818 12578
rect 2752 12268 2818 12386
rect 2752 12076 2758 12268
rect 2810 12076 2818 12268
rect 2752 11958 2818 12076
rect 2752 11766 2758 11958
rect 2810 11766 2818 11958
rect 2752 11644 2818 11766
rect 2752 11456 2758 11644
rect 2810 11456 2818 11644
rect 2752 11334 2818 11456
rect 2752 11146 2758 11334
rect 2810 11146 2818 11334
rect 2752 11026 2818 11146
rect 2752 10838 2758 11026
rect 2810 10838 2818 11026
rect 2752 10712 2818 10838
rect 2752 10526 2758 10712
rect 2810 10526 2818 10712
rect 2752 10404 2818 10526
rect 2752 10218 2758 10404
rect 2810 10218 2818 10404
rect 2752 10060 2818 10218
rect 3068 13202 3134 13358
rect 3068 13004 3074 13202
rect 3128 13004 3134 13202
rect 3068 12890 3134 13004
rect 3068 12692 3074 12890
rect 3128 12692 3134 12890
rect 3068 12578 3134 12692
rect 3068 12386 3074 12578
rect 3128 12386 3134 12578
rect 3068 12268 3134 12386
rect 3068 12076 3074 12268
rect 3126 12076 3134 12268
rect 3068 11958 3134 12076
rect 3068 11766 3074 11958
rect 3126 11766 3134 11958
rect 3068 11644 3134 11766
rect 3068 11456 3074 11644
rect 3126 11456 3134 11644
rect 3068 11334 3134 11456
rect 3068 11146 3074 11334
rect 3126 11146 3134 11334
rect 3068 11026 3134 11146
rect 3068 10838 3074 11026
rect 3126 10838 3134 11026
rect 3068 10712 3134 10838
rect 3068 10526 3074 10712
rect 3126 10526 3134 10712
rect 3068 10404 3134 10526
rect 3068 10218 3074 10404
rect 3126 10218 3134 10404
rect 3068 10060 3134 10218
rect 3384 13202 3450 13358
rect 3384 13004 3390 13202
rect 3444 13004 3450 13202
rect 3384 12890 3450 13004
rect 3384 12692 3390 12890
rect 3444 12692 3450 12890
rect 4568 12856 4662 14182
rect 69856 13822 69954 14182
rect 69866 13324 69954 13822
rect 69856 12856 69954 13324
rect 4568 12744 69954 12856
rect 3384 12578 3450 12692
rect 3384 12386 3390 12578
rect 3444 12386 3450 12578
rect 3384 12268 3450 12386
rect 3384 12076 3390 12268
rect 3442 12076 3450 12268
rect 3384 11958 3450 12076
rect 3384 11766 3390 11958
rect 3442 11766 3450 11958
rect 3384 11644 3450 11766
rect 3384 11456 3390 11644
rect 3442 11456 3450 11644
rect 3384 11334 3450 11456
rect 3384 11146 3390 11334
rect 3442 11146 3450 11334
rect 3384 11026 3450 11146
rect 3384 10838 3390 11026
rect 3442 10838 3450 11026
rect 3384 10712 3450 10838
rect 3384 10526 3390 10712
rect 3442 10526 3450 10712
rect 3384 10404 3450 10526
rect 3384 10218 3390 10404
rect 3442 10218 3450 10404
rect 3384 10060 3450 10218
rect 526 10046 3458 10060
rect 526 9994 544 10046
rect 3446 9994 3458 10046
rect 526 9982 3458 9994
rect -5724 9236 -3924 9254
rect -5724 8912 -4168 9236
rect -3986 8912 -3924 9236
rect -5724 8894 -3924 8912
rect -7574 7508 -7568 8356
rect -7368 7508 -7362 8356
rect -7574 6750 -7362 7508
rect -7574 5902 -7568 6750
rect -7368 5902 -7362 6750
rect -7574 5884 -7362 5902
rect -12170 5044 -7732 5264
rect -10226 4844 -9626 5044
rect -13830 4244 -9628 4844
rect 1750 4480 3150 9982
rect 1338 4420 3408 4480
rect 1338 4048 1370 4420
rect 1338 3740 1376 4048
rect 3362 3740 3408 4420
rect 1338 3606 3408 3740
<< via2 >>
rect -1244 31028 8992 31608
rect -17422 29110 -16842 29690
rect -16222 29110 -15642 29690
rect -15022 29110 -14442 29690
rect -13822 29110 -13242 29690
rect -12622 29110 -12042 29690
rect -11422 29110 -10842 29690
rect -10222 29110 -9642 29690
rect -9022 29110 -8442 29690
rect -7822 29110 -7242 29690
rect -6622 29110 -6042 29690
rect -5422 29110 -4842 29690
rect -18156 28872 -17580 28902
rect -18156 28472 -17786 28872
rect -17786 28472 -17590 28872
rect -17590 28472 -17580 28872
rect -18156 27960 -17580 28472
rect -18156 27266 -17580 27576
rect -18156 26866 -17786 27266
rect -17786 26866 -17590 27266
rect -17590 26866 -17580 27266
rect -18156 26554 -17580 26866
rect -18156 25660 -17580 26170
rect -18156 25260 -17786 25660
rect -17786 25260 -17590 25660
rect -17590 25260 -17580 25660
rect -18156 25148 -17580 25260
rect -18156 24054 -17580 24764
rect -18156 23742 -17786 24054
rect -17786 23742 -17590 24054
rect -17590 23742 -17580 24054
rect -18156 22448 -17580 23358
rect -18156 22336 -17786 22448
rect -17786 22336 -17590 22448
rect -17590 22336 -17580 22448
rect -18156 20930 -17580 21952
rect -18156 20442 -17786 20546
rect -17786 20442 -17590 20546
rect -17590 20442 -17580 20546
rect -18156 19524 -17580 20442
rect -18156 18836 -17786 19140
rect -17786 18836 -17590 19140
rect -17590 18836 -17580 19140
rect -18156 18118 -17580 18836
rect -18156 17630 -17580 17734
rect -18156 17230 -17786 17630
rect -17786 17230 -17590 17630
rect -17590 17230 -17580 17630
rect -18156 16712 -17580 17230
rect -18156 16024 -17580 16328
rect -18156 15624 -17786 16024
rect -17786 15624 -17590 16024
rect -17590 15624 -17580 16024
rect -18156 15306 -17580 15624
rect -18156 14418 -17580 14922
rect -18156 14018 -17786 14418
rect -17786 14018 -17590 14418
rect -17590 14018 -17580 14418
rect -18156 13900 -17580 14018
rect -16750 28872 -16174 28902
rect -16750 28472 -16380 28872
rect -16380 28472 -16184 28872
rect -16184 28472 -16174 28872
rect -16750 27960 -16174 28472
rect -16750 27266 -16174 27576
rect -16750 26866 -16380 27266
rect -16380 26866 -16184 27266
rect -16184 26866 -16174 27266
rect -16750 26554 -16174 26866
rect -16750 25660 -16174 26170
rect -16750 25260 -16380 25660
rect -16380 25260 -16184 25660
rect -16184 25260 -16174 25660
rect -16750 25148 -16174 25260
rect -16750 24054 -16174 24764
rect -16750 23742 -16380 24054
rect -16380 23742 -16184 24054
rect -16184 23742 -16174 24054
rect -16750 22448 -16174 23358
rect -16750 22336 -16380 22448
rect -16380 22336 -16184 22448
rect -16184 22336 -16174 22448
rect -16750 20930 -16174 21952
rect -16750 20442 -16380 20546
rect -16380 20442 -16184 20546
rect -16184 20442 -16174 20546
rect -16750 19524 -16174 20442
rect -16750 18836 -16380 19140
rect -16380 18836 -16184 19140
rect -16184 18836 -16174 19140
rect -16750 18118 -16174 18836
rect -16750 17630 -16174 17734
rect -16750 17230 -16380 17630
rect -16380 17230 -16184 17630
rect -16184 17230 -16174 17630
rect -16750 16712 -16174 17230
rect -16750 16024 -16174 16328
rect -16750 15624 -16380 16024
rect -16380 15624 -16184 16024
rect -16184 15624 -16174 16024
rect -16750 15306 -16174 15624
rect -16750 14418 -16174 14922
rect -16750 14018 -16380 14418
rect -16380 14018 -16184 14418
rect -16184 14018 -16174 14418
rect -16750 13900 -16174 14018
rect -15344 28872 -14768 28902
rect -15344 28472 -14974 28872
rect -14974 28472 -14778 28872
rect -14778 28472 -14768 28872
rect -15344 27960 -14768 28472
rect -15344 27266 -14768 27576
rect -15344 26866 -14974 27266
rect -14974 26866 -14778 27266
rect -14778 26866 -14768 27266
rect -15344 26554 -14768 26866
rect -15344 25660 -14768 26170
rect -15344 25260 -14974 25660
rect -14974 25260 -14778 25660
rect -14778 25260 -14768 25660
rect -15344 25148 -14768 25260
rect -15344 24054 -14768 24764
rect -15344 23742 -14974 24054
rect -14974 23742 -14778 24054
rect -14778 23742 -14768 24054
rect -15344 22448 -14768 23358
rect -15344 22336 -14974 22448
rect -14974 22336 -14778 22448
rect -14778 22336 -14768 22448
rect -15344 20930 -14768 21952
rect -15344 20442 -14974 20546
rect -14974 20442 -14778 20546
rect -14778 20442 -14768 20546
rect -15344 19524 -14768 20442
rect -15344 18836 -14974 19140
rect -14974 18836 -14778 19140
rect -14778 18836 -14768 19140
rect -15344 18118 -14768 18836
rect -15344 17630 -14768 17734
rect -15344 17230 -14974 17630
rect -14974 17230 -14778 17630
rect -14778 17230 -14768 17630
rect -15344 16712 -14768 17230
rect -15344 16024 -14768 16328
rect -15344 15624 -14974 16024
rect -14974 15624 -14778 16024
rect -14778 15624 -14768 16024
rect -15344 15306 -14768 15624
rect -15344 14418 -14768 14922
rect -15344 14018 -14974 14418
rect -14974 14018 -14778 14418
rect -14778 14018 -14768 14418
rect -15344 13900 -14768 14018
rect -13938 28872 -13362 28902
rect -13938 28472 -13568 28872
rect -13568 28472 -13372 28872
rect -13372 28472 -13362 28872
rect -13938 27960 -13362 28472
rect -13938 27266 -13362 27576
rect -13938 26866 -13568 27266
rect -13568 26866 -13372 27266
rect -13372 26866 -13362 27266
rect -13938 26554 -13362 26866
rect -13938 25660 -13362 26170
rect -13938 25260 -13568 25660
rect -13568 25260 -13372 25660
rect -13372 25260 -13362 25660
rect -13938 25148 -13362 25260
rect -13938 24054 -13362 24764
rect -13938 23742 -13568 24054
rect -13568 23742 -13372 24054
rect -13372 23742 -13362 24054
rect -13938 22448 -13362 23358
rect -13938 22336 -13568 22448
rect -13568 22336 -13372 22448
rect -13372 22336 -13362 22448
rect -13938 20930 -13362 21952
rect -13938 20442 -13568 20546
rect -13568 20442 -13372 20546
rect -13372 20442 -13362 20546
rect -13938 19524 -13362 20442
rect -13938 18836 -13568 19140
rect -13568 18836 -13372 19140
rect -13372 18836 -13362 19140
rect -13938 18118 -13362 18836
rect -13938 17630 -13362 17734
rect -13938 17230 -13568 17630
rect -13568 17230 -13372 17630
rect -13372 17230 -13362 17630
rect -13938 16712 -13362 17230
rect -13938 16024 -13362 16328
rect -13938 15624 -13568 16024
rect -13568 15624 -13372 16024
rect -13372 15624 -13362 16024
rect -13938 15306 -13362 15624
rect -13938 14418 -13362 14922
rect -13938 14018 -13568 14418
rect -13568 14018 -13372 14418
rect -13372 14018 -13362 14418
rect -13938 13900 -13362 14018
rect -12532 28872 -11956 28902
rect -12532 28472 -12162 28872
rect -12162 28472 -11966 28872
rect -11966 28472 -11956 28872
rect -12532 27960 -11956 28472
rect -12532 27266 -11956 27576
rect -12532 26866 -12162 27266
rect -12162 26866 -11966 27266
rect -11966 26866 -11956 27266
rect -12532 26554 -11956 26866
rect -12532 25660 -11956 26170
rect -12532 25260 -12162 25660
rect -12162 25260 -11966 25660
rect -11966 25260 -11956 25660
rect -12532 25148 -11956 25260
rect -12532 24054 -11956 24764
rect -12532 23742 -12162 24054
rect -12162 23742 -11966 24054
rect -11966 23742 -11956 24054
rect -12532 22448 -11956 23358
rect -12532 22336 -12162 22448
rect -12162 22336 -11966 22448
rect -11966 22336 -11956 22448
rect -12532 20930 -11956 21952
rect -12532 20442 -12162 20546
rect -12162 20442 -11966 20546
rect -11966 20442 -11956 20546
rect -12532 19524 -11956 20442
rect -12532 18836 -12162 19140
rect -12162 18836 -11966 19140
rect -11966 18836 -11956 19140
rect -12532 18118 -11956 18836
rect -12532 17630 -11956 17734
rect -12532 17230 -12162 17630
rect -12162 17230 -11966 17630
rect -11966 17230 -11956 17630
rect -12532 16712 -11956 17230
rect -12532 16024 -11956 16328
rect -12532 15624 -12162 16024
rect -12162 15624 -11966 16024
rect -11966 15624 -11956 16024
rect -12532 15306 -11956 15624
rect -12532 14418 -11956 14922
rect -12532 14018 -12162 14418
rect -12162 14018 -11966 14418
rect -11966 14018 -11956 14418
rect -12532 13900 -11956 14018
rect -11126 28872 -10550 28902
rect -11126 28472 -10756 28872
rect -10756 28472 -10560 28872
rect -10560 28472 -10550 28872
rect -11126 27960 -10550 28472
rect -11126 27266 -10550 27576
rect -11126 26866 -10756 27266
rect -10756 26866 -10560 27266
rect -10560 26866 -10550 27266
rect -11126 26554 -10550 26866
rect -11126 25660 -10550 26170
rect -11126 25260 -10756 25660
rect -10756 25260 -10560 25660
rect -10560 25260 -10550 25660
rect -11126 25148 -10550 25260
rect -11126 24054 -10550 24764
rect -11126 23742 -10756 24054
rect -10756 23742 -10560 24054
rect -10560 23742 -10550 24054
rect -11126 22448 -10550 23358
rect -11126 22336 -10756 22448
rect -10756 22336 -10560 22448
rect -10560 22336 -10550 22448
rect -11126 20930 -10550 21952
rect -11126 20442 -10756 20546
rect -10756 20442 -10560 20546
rect -10560 20442 -10550 20546
rect -11126 19524 -10550 20442
rect -11126 18836 -10756 19140
rect -10756 18836 -10560 19140
rect -10560 18836 -10550 19140
rect -11126 18118 -10550 18836
rect -11126 17630 -10550 17734
rect -11126 17230 -10756 17630
rect -10756 17230 -10560 17630
rect -10560 17230 -10550 17630
rect -11126 16712 -10550 17230
rect -11126 16024 -10550 16328
rect -11126 15624 -10756 16024
rect -10756 15624 -10560 16024
rect -10560 15624 -10550 16024
rect -11126 15306 -10550 15624
rect -11126 14418 -10550 14922
rect -11126 14018 -10756 14418
rect -10756 14018 -10560 14418
rect -10560 14018 -10550 14418
rect -11126 13900 -10550 14018
rect -9720 28872 -9144 28902
rect -9720 28472 -9350 28872
rect -9350 28472 -9154 28872
rect -9154 28472 -9144 28872
rect -9720 27960 -9144 28472
rect -9720 27266 -9144 27576
rect -9720 26866 -9350 27266
rect -9350 26866 -9154 27266
rect -9154 26866 -9144 27266
rect -9720 26554 -9144 26866
rect -9720 25660 -9144 26170
rect -9720 25260 -9350 25660
rect -9350 25260 -9154 25660
rect -9154 25260 -9144 25660
rect -9720 25148 -9144 25260
rect -9720 24054 -9144 24764
rect -9720 23742 -9350 24054
rect -9350 23742 -9154 24054
rect -9154 23742 -9144 24054
rect -9720 22448 -9144 23358
rect -9720 22336 -9350 22448
rect -9350 22336 -9154 22448
rect -9154 22336 -9144 22448
rect -9720 20930 -9144 21952
rect -9720 20442 -9350 20546
rect -9350 20442 -9154 20546
rect -9154 20442 -9144 20546
rect -9720 19524 -9144 20442
rect -9720 18836 -9350 19140
rect -9350 18836 -9154 19140
rect -9154 18836 -9144 19140
rect -9720 18118 -9144 18836
rect -9720 17630 -9144 17734
rect -9720 17230 -9350 17630
rect -9350 17230 -9154 17630
rect -9154 17230 -9144 17630
rect -9720 16712 -9144 17230
rect -9720 16024 -9144 16328
rect -9720 15624 -9350 16024
rect -9350 15624 -9154 16024
rect -9154 15624 -9144 16024
rect -9720 15306 -9144 15624
rect -9720 14418 -9144 14922
rect -9720 14018 -9350 14418
rect -9350 14018 -9154 14418
rect -9154 14018 -9144 14418
rect -9720 13900 -9144 14018
rect -8314 28872 -7738 28902
rect -8314 28472 -7944 28872
rect -7944 28472 -7748 28872
rect -7748 28472 -7738 28872
rect -8314 27960 -7738 28472
rect -8314 27266 -7738 27576
rect -8314 26866 -7944 27266
rect -7944 26866 -7748 27266
rect -7748 26866 -7738 27266
rect -8314 26554 -7738 26866
rect -8314 25660 -7738 26170
rect -8314 25260 -7944 25660
rect -7944 25260 -7748 25660
rect -7748 25260 -7738 25660
rect -8314 25148 -7738 25260
rect -8314 24054 -7738 24764
rect -8314 23742 -7944 24054
rect -7944 23742 -7748 24054
rect -7748 23742 -7738 24054
rect -8314 22448 -7738 23358
rect -8314 22336 -7944 22448
rect -7944 22336 -7748 22448
rect -7748 22336 -7738 22448
rect -8314 20930 -7738 21952
rect -8314 20442 -7944 20546
rect -7944 20442 -7748 20546
rect -7748 20442 -7738 20546
rect -8314 19524 -7738 20442
rect -8314 18836 -7944 19140
rect -7944 18836 -7748 19140
rect -7748 18836 -7738 19140
rect -8314 18118 -7738 18836
rect -8314 17630 -7738 17734
rect -8314 17230 -7944 17630
rect -7944 17230 -7748 17630
rect -7748 17230 -7738 17630
rect -8314 16712 -7738 17230
rect -8314 16024 -7738 16328
rect -8314 15624 -7944 16024
rect -7944 15624 -7748 16024
rect -7748 15624 -7738 16024
rect -8314 15306 -7738 15624
rect -8314 14418 -7738 14922
rect -8314 14018 -7944 14418
rect -7944 14018 -7748 14418
rect -7748 14018 -7738 14418
rect -8314 13900 -7738 14018
rect -6908 28872 -6332 28902
rect -6908 28472 -6538 28872
rect -6538 28472 -6342 28872
rect -6342 28472 -6332 28872
rect -6908 27960 -6332 28472
rect -6908 27266 -6332 27576
rect -6908 26866 -6538 27266
rect -6538 26866 -6342 27266
rect -6342 26866 -6332 27266
rect -6908 26554 -6332 26866
rect -6908 25660 -6332 26170
rect -6908 25260 -6538 25660
rect -6538 25260 -6342 25660
rect -6342 25260 -6332 25660
rect -6908 25148 -6332 25260
rect -6908 24054 -6332 24764
rect -6908 23742 -6538 24054
rect -6538 23742 -6342 24054
rect -6342 23742 -6332 24054
rect -6908 22448 -6332 23358
rect -6908 22336 -6538 22448
rect -6538 22336 -6342 22448
rect -6342 22336 -6332 22448
rect -6908 20930 -6332 21952
rect -6908 20442 -6538 20546
rect -6538 20442 -6342 20546
rect -6342 20442 -6332 20546
rect -6908 19524 -6332 20442
rect -6908 18836 -6538 19140
rect -6538 18836 -6342 19140
rect -6342 18836 -6332 19140
rect -6908 18118 -6332 18836
rect -6908 17630 -6332 17734
rect -6908 17230 -6538 17630
rect -6538 17230 -6342 17630
rect -6342 17230 -6332 17630
rect -6908 16712 -6332 17230
rect -6908 16024 -6332 16328
rect -6908 15624 -6538 16024
rect -6538 15624 -6342 16024
rect -6342 15624 -6332 16024
rect -6908 15306 -6332 15624
rect -6908 14418 -6332 14922
rect -6908 14018 -6538 14418
rect -6538 14018 -6342 14418
rect -6342 14018 -6332 14418
rect -6908 13900 -6332 14018
rect -5502 28872 -4926 28902
rect -5502 28472 -5132 28872
rect -5132 28472 -4936 28872
rect -4936 28472 -4926 28872
rect -5502 27960 -4926 28472
rect -5502 27266 -4926 27576
rect -5502 26866 -5132 27266
rect -5132 26866 -4936 27266
rect -4936 26866 -4926 27266
rect -5502 26554 -4926 26866
rect -5502 25660 -4926 26170
rect -5502 25260 -5132 25660
rect -5132 25260 -4936 25660
rect -4936 25260 -4926 25660
rect -5502 25148 -4926 25260
rect -5502 24054 -4926 24764
rect -5502 23742 -5132 24054
rect -5132 23742 -4936 24054
rect -4936 23742 -4926 24054
rect -5502 22448 -4926 23358
rect -5502 22336 -5132 22448
rect -5132 22336 -4936 22448
rect -4936 22336 -4926 22448
rect -5502 20930 -4926 21952
rect -5502 20442 -5132 20546
rect -5132 20442 -4936 20546
rect -4936 20442 -4926 20546
rect -5502 19524 -4926 20442
rect -5502 18836 -5132 19140
rect -5132 18836 -4936 19140
rect -4936 18836 -4926 19140
rect -5502 18118 -4926 18836
rect -5502 17630 -4926 17734
rect -5502 17230 -5132 17630
rect -5132 17230 -4936 17630
rect -4936 17230 -4926 17630
rect -5502 16712 -4926 17230
rect -5502 16024 -4926 16328
rect -5502 15624 -5132 16024
rect -5132 15624 -4936 16024
rect -4936 15624 -4926 16024
rect -5502 15306 -4926 15624
rect -5502 14418 -4926 14922
rect -5502 14018 -5132 14418
rect -5132 14018 -4936 14418
rect -4936 14018 -4926 14418
rect -5502 13900 -4926 14018
rect -3870 28490 -3290 29690
rect -17826 13202 -17226 13206
rect -16826 13202 -16160 13206
rect -15826 13202 -14226 13206
rect -13948 13202 -13226 13206
rect -12826 13202 -11942 13206
rect -11826 13202 -11226 13206
rect -11136 13202 -10226 13206
rect -9826 13202 -9130 13206
rect -8826 13202 -7226 13206
rect -6918 13202 -6226 13206
rect -5826 13202 -4912 13206
rect -18156 12606 -4912 13202
rect -2982 24656 -2396 30034
rect -1224 29300 -444 30080
rect 172 29300 952 30080
rect 1568 29300 2348 30080
rect 2964 29300 3744 30080
rect -1696 28878 -1368 29106
rect -300 28878 28 29106
rect 1096 28878 1424 29106
rect 2492 28878 2820 29106
rect 3888 28878 4216 29106
rect -1224 27904 -444 28684
rect 172 27904 952 28684
rect 1568 27904 2348 28684
rect 2964 27904 3744 28684
rect -1696 27482 -1368 27710
rect -300 27482 28 27710
rect 1096 27482 1424 27710
rect 2492 27482 2820 27710
rect 3888 27482 4216 27710
rect -1224 26508 -444 27288
rect 172 26508 952 27288
rect 1568 26508 2348 27288
rect 2964 26508 3744 27288
rect 8992 28728 50182 29308
rect 9920 28122 10500 28166
rect 9920 27342 10500 28122
rect 9920 26726 10500 27342
rect -1696 26086 -1368 26314
rect -300 26086 28 26314
rect 1096 26086 1424 26314
rect 2492 26086 2820 26314
rect 3888 26086 4216 26314
rect -1224 25112 -444 25892
rect 172 25112 952 25892
rect 1568 25112 2348 25892
rect 2964 25112 3744 25892
rect 9920 25946 10500 26726
rect -1696 24690 -1368 24918
rect -300 24690 28 24918
rect 1096 24690 1424 24918
rect 2492 24690 2820 24918
rect 3888 24690 4216 24918
rect 9920 24774 10500 25946
rect 10796 25716 11020 28256
rect 11316 28122 11896 28166
rect 11316 27342 11896 28122
rect 11316 26726 11896 27342
rect 11316 25946 11896 26726
rect 11316 24774 11896 25946
rect 12192 25716 12416 28256
rect 12712 28122 13292 28166
rect 12712 27342 13292 28122
rect 12712 26726 13292 27342
rect 12712 25946 13292 26726
rect 12712 24774 13292 25946
rect 13588 25716 13812 28256
rect 14108 28122 14688 28166
rect 14108 27342 14688 28122
rect 14108 26726 14688 27342
rect 14108 25946 14688 26726
rect 14108 24774 14688 25946
rect 14984 25716 15208 28256
rect 15504 28122 16084 28166
rect 15504 27342 16084 28122
rect 15504 26726 16084 27342
rect 15504 25946 16084 26726
rect 15504 24774 16084 25946
rect 16380 25716 16604 28256
rect 16900 28122 17480 28166
rect 16900 27342 17480 28122
rect 16900 26726 17480 27342
rect 16900 25946 17480 26726
rect 16900 24774 17480 25946
rect 17776 25716 18000 28256
rect 18296 28122 18876 28166
rect 18296 27342 18876 28122
rect 18296 26726 18876 27342
rect 18296 25946 18876 26726
rect 18296 24774 18876 25946
rect 19172 25716 19396 28256
rect 19692 28122 20272 28166
rect 19692 27342 20272 28122
rect 19692 26726 20272 27342
rect 19692 25946 20272 26726
rect 19692 24774 20272 25946
rect 20568 25716 20792 28256
rect 21088 28122 21668 28166
rect 21088 27342 21668 28122
rect 21088 26726 21668 27342
rect 21088 25946 21668 26726
rect 21088 24774 21668 25946
rect 21964 25716 22188 28256
rect 22484 28122 23064 28166
rect 22484 27342 23064 28122
rect 22484 26726 23064 27342
rect 22484 25946 23064 26726
rect 22484 24774 23064 25946
rect 23360 25716 23584 28256
rect 23880 28122 24460 28166
rect 23880 27342 24460 28122
rect 23880 26726 24460 27342
rect 23880 25946 24460 26726
rect 23880 24774 24460 25946
rect 24756 25716 24980 28256
rect 25276 28122 25856 28166
rect 25276 27342 25856 28122
rect 25276 26726 25856 27342
rect 25276 25946 25856 26726
rect 25276 24774 25856 25946
rect 26152 25716 26376 28256
rect 26672 28122 27252 28166
rect 26672 27342 27252 28122
rect 26672 26726 27252 27342
rect 26672 25946 27252 26726
rect 26672 24774 27252 25946
rect 27548 25716 27772 28256
rect 28068 28122 28648 28166
rect 28068 27342 28648 28122
rect 28068 26726 28648 27342
rect 28068 25946 28648 26726
rect 28068 24774 28648 25946
rect 28944 25716 29168 28256
rect 29464 28122 30044 28166
rect 29464 27342 30044 28122
rect 29464 26726 30044 27342
rect 29464 25946 30044 26726
rect 29464 24774 30044 25946
rect 30340 25716 30564 28256
rect 30860 28122 31440 28166
rect 30860 27342 31440 28122
rect 30860 26726 31440 27342
rect 30860 25946 31440 26726
rect 30860 24774 31440 25946
rect 31736 25716 31960 28256
rect 32256 28122 32836 28166
rect 32256 27342 32836 28122
rect 32256 26726 32836 27342
rect 32256 25946 32836 26726
rect 32256 24774 32836 25946
rect 33132 25716 33356 28256
rect 33652 28122 34232 28166
rect 33652 27342 34232 28122
rect 33652 26726 34232 27342
rect 33652 25946 34232 26726
rect 33652 24774 34232 25946
rect 34528 25716 34752 28256
rect 35048 28122 35628 28166
rect 35048 27342 35628 28122
rect 35048 26726 35628 27342
rect 35048 25946 35628 26726
rect 35048 24774 35628 25946
rect 35924 25716 36148 28256
rect 36444 28122 37024 28166
rect 36444 27342 37024 28122
rect 36444 26726 37024 27342
rect 36444 25946 37024 26726
rect 36444 24774 37024 25946
rect 37320 25716 37544 28256
rect 37840 28122 38420 28166
rect 37840 27342 38420 28122
rect 37840 26726 38420 27342
rect 37840 25946 38420 26726
rect 37840 24774 38420 25946
rect 38716 25716 38940 28256
rect 39236 28122 39816 28166
rect 39236 27342 39816 28122
rect 39236 26726 39816 27342
rect 39236 25946 39816 26726
rect 39236 24774 39816 25946
rect 40112 25716 40336 28256
rect 40632 28122 41212 28166
rect 40632 27342 41212 28122
rect 40632 26726 41212 27342
rect 40632 25946 41212 26726
rect 40632 24774 41212 25946
rect 41508 25716 41732 28256
rect 42028 28122 42608 28166
rect 42028 27342 42608 28122
rect 42028 26726 42608 27342
rect 42028 25946 42608 26726
rect 42028 24774 42608 25946
rect 42904 25716 43128 28256
rect 43424 28122 44004 28166
rect 43424 27342 44004 28122
rect 43424 26726 44004 27342
rect 43424 25946 44004 26726
rect 43424 24774 44004 25946
rect 44300 25716 44524 28256
rect 44820 28122 45400 28166
rect 44820 27342 45400 28122
rect 44820 26726 45400 27342
rect 44820 25946 45400 26726
rect 44820 24774 45400 25946
rect 45696 25716 45920 28256
rect 46216 28122 46796 28166
rect 46216 27342 46796 28122
rect 46216 26726 46796 27342
rect 46216 25946 46796 26726
rect 46216 24774 46796 25946
rect 47092 25716 47316 28256
rect 47612 28122 48192 28166
rect 47612 27342 48192 28122
rect 47612 26726 48192 27342
rect 47612 25946 48192 26726
rect 47612 24774 48192 25946
rect 48488 25716 48712 28256
rect 49008 28122 49588 28166
rect 49008 27342 49588 28122
rect 49008 26726 49588 27342
rect 49008 25946 49588 26726
rect 49008 24774 49588 25946
rect 49884 25716 50108 28256
rect 50404 28122 50984 28166
rect 50404 27342 50984 28122
rect 50404 26726 50984 27342
rect 50404 25946 50984 26726
rect 50404 24774 50984 25946
rect -1228 23856 3618 24438
rect 4642 24394 70084 24774
rect 3703 22941 4093 23331
rect -2963 18645 -2573 19035
rect -3870 11686 -3290 12886
rect 4662 13822 69856 14182
rect 4662 13324 69410 13822
rect 69410 13324 69856 13822
rect 4662 12856 69856 13324
rect 1370 4048 3362 4420
rect 1376 3740 3362 4048
<< metal3 >>
rect -1254 31608 9582 31618
rect -1254 31028 -1244 31608
rect 8992 31028 9582 31608
rect -1254 31018 9582 31028
rect 3928 30186 4298 31018
rect 4586 30186 5186 31018
rect -1234 30080 -434 30090
rect -2992 30034 -2386 30044
rect -17432 29690 -3280 29700
rect -17432 29110 -17422 29690
rect -16842 29110 -16222 29690
rect -15642 29110 -15022 29690
rect -14442 29110 -13822 29690
rect -13242 29110 -12622 29690
rect -12042 29110 -11422 29690
rect -10842 29110 -10222 29690
rect -9642 29110 -9022 29690
rect -8442 29110 -7822 29690
rect -7242 29110 -6622 29690
rect -6042 29110 -5422 29690
rect -4842 29110 -3870 29690
rect -17432 29100 -3870 29110
rect -18166 28902 -17566 28910
rect -18166 27960 -18156 28902
rect -17580 27960 -17566 28902
rect -18166 27576 -17566 27960
rect -18166 26554 -18156 27576
rect -17580 26554 -17566 27576
rect -18166 26170 -17566 26554
rect -18166 25148 -18156 26170
rect -17580 25148 -17566 26170
rect -18166 24764 -17566 25148
rect -18166 23742 -18156 24764
rect -17580 23742 -17566 24764
rect -18166 23358 -17566 23742
rect -18166 22336 -18156 23358
rect -17580 22336 -17566 23358
rect -18166 21952 -17566 22336
rect -18166 20930 -18156 21952
rect -17580 20930 -17566 21952
rect -18166 20546 -17566 20930
rect -18166 19524 -18156 20546
rect -17580 19524 -17566 20546
rect -18166 19140 -17566 19524
rect -18166 18118 -18156 19140
rect -17580 18118 -17566 19140
rect -18166 17734 -17566 18118
rect -18166 16712 -18156 17734
rect -17580 16712 -17566 17734
rect -18166 16328 -17566 16712
rect -18166 15306 -18156 16328
rect -17580 15306 -17566 16328
rect -18166 14922 -17566 15306
rect -18166 13900 -18156 14922
rect -17580 13900 -17566 14922
rect -18166 13212 -17566 13900
rect -16760 28902 -16160 28910
rect -16760 27960 -16750 28902
rect -16174 27960 -16160 28902
rect -16760 27576 -16160 27960
rect -16760 26554 -16750 27576
rect -16174 26554 -16160 27576
rect -16760 26170 -16160 26554
rect -16760 25148 -16750 26170
rect -16174 25148 -16160 26170
rect -16760 24764 -16160 25148
rect -16760 23742 -16750 24764
rect -16174 23742 -16160 24764
rect -16760 23358 -16160 23742
rect -16760 22336 -16750 23358
rect -16174 22336 -16160 23358
rect -16760 21952 -16160 22336
rect -16760 20930 -16750 21952
rect -16174 20930 -16160 21952
rect -16760 20546 -16160 20930
rect -16760 19524 -16750 20546
rect -16174 19524 -16160 20546
rect -16760 19140 -16160 19524
rect -16760 18118 -16750 19140
rect -16174 18118 -16160 19140
rect -16760 17734 -16160 18118
rect -16760 16712 -16750 17734
rect -16174 16712 -16160 17734
rect -16760 16328 -16160 16712
rect -16760 15306 -16750 16328
rect -16174 15306 -16160 16328
rect -16760 14922 -16160 15306
rect -16760 13900 -16750 14922
rect -16174 13900 -16160 14922
rect -16760 13212 -16160 13900
rect -15354 28902 -14754 28910
rect -15354 27960 -15344 28902
rect -14768 27960 -14754 28902
rect -15354 27576 -14754 27960
rect -15354 26554 -15344 27576
rect -14768 26554 -14754 27576
rect -15354 26170 -14754 26554
rect -15354 25148 -15344 26170
rect -14768 25148 -14754 26170
rect -15354 24764 -14754 25148
rect -15354 23742 -15344 24764
rect -14768 23742 -14754 24764
rect -15354 23358 -14754 23742
rect -15354 22336 -15344 23358
rect -14768 22336 -14754 23358
rect -15354 21952 -14754 22336
rect -15354 20930 -15344 21952
rect -14768 20930 -14754 21952
rect -15354 20546 -14754 20930
rect -15354 19524 -15344 20546
rect -14768 19524 -14754 20546
rect -15354 19140 -14754 19524
rect -15354 18118 -15344 19140
rect -14768 18118 -14754 19140
rect -15354 17734 -14754 18118
rect -15354 16712 -15344 17734
rect -14768 16712 -14754 17734
rect -15354 16328 -14754 16712
rect -15354 15306 -15344 16328
rect -14768 15306 -14754 16328
rect -15354 14922 -14754 15306
rect -15354 13900 -15344 14922
rect -14768 13900 -14754 14922
rect -15354 13212 -14754 13900
rect -13948 28902 -13348 28910
rect -13948 27960 -13938 28902
rect -13362 27960 -13348 28902
rect -13948 27576 -13348 27960
rect -13948 26554 -13938 27576
rect -13362 26554 -13348 27576
rect -13948 26170 -13348 26554
rect -13948 25148 -13938 26170
rect -13362 25148 -13348 26170
rect -13948 24764 -13348 25148
rect -13948 23742 -13938 24764
rect -13362 23742 -13348 24764
rect -13948 23358 -13348 23742
rect -13948 22336 -13938 23358
rect -13362 22336 -13348 23358
rect -13948 21952 -13348 22336
rect -13948 20930 -13938 21952
rect -13362 20930 -13348 21952
rect -13948 20546 -13348 20930
rect -13948 19524 -13938 20546
rect -13362 19524 -13348 20546
rect -13948 19140 -13348 19524
rect -13948 18118 -13938 19140
rect -13362 18118 -13348 19140
rect -13948 17734 -13348 18118
rect -13948 16712 -13938 17734
rect -13362 16712 -13348 17734
rect -13948 16328 -13348 16712
rect -13948 15306 -13938 16328
rect -13362 15306 -13348 16328
rect -13948 14922 -13348 15306
rect -13948 13900 -13938 14922
rect -13362 13900 -13348 14922
rect -13948 13212 -13348 13900
rect -12542 28902 -11942 28910
rect -12542 27960 -12532 28902
rect -11956 27960 -11942 28902
rect -12542 27576 -11942 27960
rect -12542 26554 -12532 27576
rect -11956 26554 -11942 27576
rect -12542 26170 -11942 26554
rect -12542 25148 -12532 26170
rect -11956 25148 -11942 26170
rect -12542 24764 -11942 25148
rect -12542 23742 -12532 24764
rect -11956 23742 -11942 24764
rect -12542 23358 -11942 23742
rect -12542 22336 -12532 23358
rect -11956 22336 -11942 23358
rect -12542 21952 -11942 22336
rect -12542 20930 -12532 21952
rect -11956 20930 -11942 21952
rect -12542 20546 -11942 20930
rect -12542 19524 -12532 20546
rect -11956 19524 -11942 20546
rect -12542 19140 -11942 19524
rect -12542 18118 -12532 19140
rect -11956 18118 -11942 19140
rect -12542 17734 -11942 18118
rect -12542 16712 -12532 17734
rect -11956 16712 -11942 17734
rect -12542 16328 -11942 16712
rect -12542 15306 -12532 16328
rect -11956 15306 -11942 16328
rect -12542 14922 -11942 15306
rect -12542 13900 -12532 14922
rect -11956 13900 -11942 14922
rect -12542 13212 -11942 13900
rect -11136 28902 -10536 28910
rect -11136 27960 -11126 28902
rect -10550 27960 -10536 28902
rect -11136 27576 -10536 27960
rect -11136 26554 -11126 27576
rect -10550 26554 -10536 27576
rect -11136 26170 -10536 26554
rect -11136 25148 -11126 26170
rect -10550 25148 -10536 26170
rect -11136 24764 -10536 25148
rect -11136 23742 -11126 24764
rect -10550 23742 -10536 24764
rect -11136 23358 -10536 23742
rect -11136 22336 -11126 23358
rect -10550 22336 -10536 23358
rect -11136 21952 -10536 22336
rect -11136 20930 -11126 21952
rect -10550 20930 -10536 21952
rect -11136 20546 -10536 20930
rect -11136 19524 -11126 20546
rect -10550 19524 -10536 20546
rect -11136 19140 -10536 19524
rect -11136 18118 -11126 19140
rect -10550 18118 -10536 19140
rect -11136 17734 -10536 18118
rect -11136 16712 -11126 17734
rect -10550 16712 -10536 17734
rect -11136 16328 -10536 16712
rect -11136 15306 -11126 16328
rect -10550 15306 -10536 16328
rect -11136 14922 -10536 15306
rect -11136 13900 -11126 14922
rect -10550 13900 -10536 14922
rect -11136 13212 -10536 13900
rect -9730 28902 -9130 28910
rect -9730 27960 -9720 28902
rect -9144 27960 -9130 28902
rect -9730 27576 -9130 27960
rect -9730 26554 -9720 27576
rect -9144 26554 -9130 27576
rect -9730 26170 -9130 26554
rect -9730 25148 -9720 26170
rect -9144 25148 -9130 26170
rect -9730 24764 -9130 25148
rect -9730 23742 -9720 24764
rect -9144 23742 -9130 24764
rect -9730 23358 -9130 23742
rect -9730 22336 -9720 23358
rect -9144 22336 -9130 23358
rect -9730 21952 -9130 22336
rect -9730 20930 -9720 21952
rect -9144 20930 -9130 21952
rect -9730 20546 -9130 20930
rect -9730 19524 -9720 20546
rect -9144 19524 -9130 20546
rect -9730 19140 -9130 19524
rect -9730 18118 -9720 19140
rect -9144 18118 -9130 19140
rect -9730 17734 -9130 18118
rect -9730 16712 -9720 17734
rect -9144 16712 -9130 17734
rect -9730 16328 -9130 16712
rect -9730 15306 -9720 16328
rect -9144 15306 -9130 16328
rect -9730 14922 -9130 15306
rect -9730 13900 -9720 14922
rect -9144 13900 -9130 14922
rect -9730 13212 -9130 13900
rect -8324 28902 -7724 28910
rect -8324 27960 -8314 28902
rect -7738 27960 -7724 28902
rect -8324 27576 -7724 27960
rect -8324 26554 -8314 27576
rect -7738 26554 -7724 27576
rect -8324 26170 -7724 26554
rect -8324 25148 -8314 26170
rect -7738 25148 -7724 26170
rect -8324 24764 -7724 25148
rect -8324 23742 -8314 24764
rect -7738 23742 -7724 24764
rect -8324 23358 -7724 23742
rect -8324 22336 -8314 23358
rect -7738 22336 -7724 23358
rect -8324 21952 -7724 22336
rect -8324 20930 -8314 21952
rect -7738 20930 -7724 21952
rect -8324 20546 -7724 20930
rect -8324 19524 -8314 20546
rect -7738 19524 -7724 20546
rect -8324 19140 -7724 19524
rect -8324 18118 -8314 19140
rect -7738 18118 -7724 19140
rect -8324 17734 -7724 18118
rect -8324 16712 -8314 17734
rect -7738 16712 -7724 17734
rect -8324 16328 -7724 16712
rect -8324 15306 -8314 16328
rect -7738 15306 -7724 16328
rect -8324 14922 -7724 15306
rect -8324 13900 -8314 14922
rect -7738 13900 -7724 14922
rect -8324 13212 -7724 13900
rect -6918 28902 -6318 28910
rect -6918 27960 -6908 28902
rect -6332 27960 -6318 28902
rect -6918 27576 -6318 27960
rect -6918 26554 -6908 27576
rect -6332 26554 -6318 27576
rect -6918 26170 -6318 26554
rect -6918 25148 -6908 26170
rect -6332 25148 -6318 26170
rect -6918 24764 -6318 25148
rect -6918 23742 -6908 24764
rect -6332 23742 -6318 24764
rect -6918 23358 -6318 23742
rect -6918 22336 -6908 23358
rect -6332 22336 -6318 23358
rect -6918 21952 -6318 22336
rect -6918 20930 -6908 21952
rect -6332 20930 -6318 21952
rect -6918 20546 -6318 20930
rect -6918 19524 -6908 20546
rect -6332 19524 -6318 20546
rect -6918 19140 -6318 19524
rect -6918 18118 -6908 19140
rect -6332 18118 -6318 19140
rect -6918 17734 -6318 18118
rect -6918 16712 -6908 17734
rect -6332 16712 -6318 17734
rect -6918 16328 -6318 16712
rect -6918 15306 -6908 16328
rect -6332 15306 -6318 16328
rect -6918 14922 -6318 15306
rect -6918 13900 -6908 14922
rect -6332 13900 -6318 14922
rect -6918 13212 -6318 13900
rect -5512 28902 -4912 28910
rect -5512 27960 -5502 28902
rect -4926 27960 -4912 28902
rect -5512 27576 -4912 27960
rect -5512 26554 -5502 27576
rect -4926 26554 -4912 27576
rect -5512 26170 -4912 26554
rect -5512 25148 -5502 26170
rect -4926 25148 -4912 26170
rect -5512 24764 -4912 25148
rect -5512 23742 -5502 24764
rect -4926 23742 -4912 24764
rect -5512 23358 -4912 23742
rect -5512 22336 -5502 23358
rect -4926 22336 -4912 23358
rect -5512 21952 -4912 22336
rect -5512 20930 -5502 21952
rect -4926 20930 -4912 21952
rect -5512 20546 -4912 20930
rect -5512 19524 -5502 20546
rect -4926 19524 -4912 20546
rect -5512 19140 -4912 19524
rect -5512 18118 -5502 19140
rect -4926 18118 -4912 19140
rect -5512 17734 -4912 18118
rect -5512 16712 -5502 17734
rect -4926 16712 -4912 17734
rect -5512 16328 -4912 16712
rect -5512 15306 -5502 16328
rect -4926 15306 -4912 16328
rect -5512 14922 -4912 15306
rect -5512 13900 -5502 14922
rect -4926 13900 -4912 14922
rect -5512 13216 -4912 13900
rect -3880 28490 -3870 29100
rect -3290 28490 -3280 29690
rect -5512 13212 -4900 13216
rect -18166 13206 -4900 13212
rect -18166 13202 -17826 13206
rect -17226 13202 -16826 13206
rect -16160 13202 -15826 13206
rect -14226 13202 -13948 13206
rect -13226 13202 -12826 13206
rect -11942 13202 -11826 13206
rect -11226 13202 -11136 13206
rect -10226 13202 -9826 13206
rect -9130 13202 -8826 13206
rect -7226 13202 -6918 13206
rect -6226 13202 -5826 13206
rect -18166 12606 -18156 13202
rect -4912 12606 -4900 13206
rect -18166 12596 -4900 12606
rect -3880 12886 -3280 28490
rect -2992 24656 -2982 30034
rect -2396 29990 -2386 30034
rect -1234 29990 -1224 30080
rect -2396 29390 -1224 29990
rect -2396 28594 -2386 29390
rect -1234 29300 -1224 29390
rect -444 29990 -434 30080
rect 162 30080 962 30090
rect 162 29990 172 30080
rect -444 29390 172 29990
rect -444 29300 -434 29390
rect -1234 29290 -434 29300
rect 162 29300 172 29390
rect 952 29990 962 30080
rect 1558 30080 2358 30090
rect 1558 29990 1568 30080
rect 952 29390 1568 29990
rect 952 29300 962 29390
rect 162 29290 962 29300
rect 1558 29300 1568 29390
rect 2348 29990 2358 30080
rect 2954 30080 3754 30090
rect 2954 29990 2964 30080
rect 2348 29390 2964 29990
rect 2348 29300 2358 29390
rect 1558 29290 2358 29300
rect 2954 29300 2964 29390
rect 3744 29300 3754 30080
rect 2954 29290 3754 29300
rect 3928 29586 5186 30186
rect 3928 29386 4298 29586
rect 5384 29386 5984 31018
rect 3928 29116 5984 29386
rect -1780 29106 5984 29116
rect -1780 28878 -1696 29106
rect -1368 28878 -300 29106
rect 28 28878 1096 29106
rect 1424 28878 2492 29106
rect 2820 28878 3888 29106
rect 4216 28878 5984 29106
rect -1780 28868 5984 28878
rect 3928 28786 5984 28868
rect -1234 28684 -434 28694
rect -1234 28594 -1224 28684
rect -2396 27994 -1224 28594
rect -2396 27198 -2386 27994
rect -1234 27904 -1224 27994
rect -444 28594 -434 28684
rect 162 28684 962 28694
rect 162 28594 172 28684
rect -444 27994 172 28594
rect -444 27904 -434 27994
rect -1234 27894 -434 27904
rect 162 27904 172 27994
rect 952 28594 962 28684
rect 1558 28684 2358 28694
rect 1558 28594 1568 28684
rect 952 27994 1568 28594
rect 952 27904 962 27994
rect 162 27894 962 27904
rect 1558 27904 1568 27994
rect 2348 28594 2358 28684
rect 2954 28684 3754 28694
rect 2954 28594 2964 28684
rect 2348 27994 2964 28594
rect 2348 27904 2358 27994
rect 1558 27894 2358 27904
rect 2954 27904 2964 27994
rect 3744 27904 3754 28684
rect 2954 27894 3754 27904
rect 3928 28586 4298 28786
rect 5384 28784 5984 28786
rect 6184 28586 6784 31018
rect 3928 27986 6784 28586
rect 3928 27786 4298 27986
rect 6184 27984 6784 27986
rect 6984 27786 7584 31018
rect 3928 27720 7584 27786
rect -1780 27710 7584 27720
rect -1780 27482 -1696 27710
rect -1368 27482 -300 27710
rect 28 27482 1096 27710
rect 1424 27482 2492 27710
rect 2820 27482 3888 27710
rect 4216 27482 7584 27710
rect -1780 27472 7584 27482
rect -1234 27288 -434 27298
rect -1234 27198 -1224 27288
rect -2396 26598 -1224 27198
rect -2396 25802 -2386 26598
rect -1234 26508 -1224 26598
rect -444 27198 -434 27288
rect 162 27288 962 27298
rect 162 27198 172 27288
rect -444 26598 172 27198
rect -444 26508 -434 26598
rect -1234 26498 -434 26508
rect 162 26508 172 26598
rect 952 27198 962 27288
rect 1558 27288 2358 27298
rect 1558 27198 1568 27288
rect 952 26598 1568 27198
rect 952 26508 962 26598
rect 162 26498 962 26508
rect 1558 26508 1568 26598
rect 2348 27198 2358 27288
rect 2954 27288 3754 27298
rect 2954 27198 2964 27288
rect 2348 26598 2964 27198
rect 2348 26508 2358 26598
rect 1558 26498 2358 26508
rect 2954 26508 2964 26598
rect 3744 26508 3754 27288
rect 2954 26498 3754 26508
rect 3928 27186 7584 27472
rect 3928 26986 4298 27186
rect 6984 27184 7584 27186
rect 7784 26986 8384 31018
rect 8982 29318 9582 31018
rect 8982 29308 50192 29318
rect 8982 28728 8992 29308
rect 50182 28728 50192 29308
rect 8982 28718 50192 28728
rect 10784 28256 11032 28718
rect 3928 26386 8384 26986
rect 3928 26324 4298 26386
rect 7784 26384 8384 26386
rect 9910 28166 10510 28176
rect -1780 26314 4298 26324
rect -1780 26086 -1696 26314
rect -1368 26086 -300 26314
rect 28 26086 1096 26314
rect 1424 26086 2492 26314
rect 2820 26086 3888 26314
rect 4216 26086 4298 26314
rect -1780 26076 4298 26086
rect -1234 25892 -434 25902
rect -1234 25802 -1224 25892
rect -2396 25202 -1224 25802
rect -2396 24656 -2386 25202
rect -1234 25112 -1224 25202
rect -444 25802 -434 25892
rect 162 25892 962 25902
rect 162 25802 172 25892
rect -444 25202 172 25802
rect -444 25112 -434 25202
rect -1234 25102 -434 25112
rect 162 25112 172 25202
rect 952 25802 962 25892
rect 1558 25892 2358 25902
rect 1558 25802 1568 25892
rect 952 25202 1568 25802
rect 952 25112 962 25202
rect 162 25102 962 25112
rect 1558 25112 1568 25202
rect 2348 25802 2358 25892
rect 2954 25892 3754 25902
rect 2954 25802 2964 25892
rect 2348 25202 2964 25802
rect 2348 25112 2358 25202
rect 1558 25102 2358 25112
rect 2954 25112 2964 25202
rect 3744 25112 3754 25892
rect 2954 25102 3754 25112
rect 3928 24928 4298 26076
rect -2992 24446 -2386 24656
rect -1780 24918 4298 24928
rect -1780 24690 -1696 24918
rect -1368 24690 -300 24918
rect 28 24690 1096 24918
rect 1424 24690 2492 24918
rect 2820 24690 3888 24918
rect 4216 24690 4298 24918
rect 9910 24784 9920 28166
rect -1780 24556 4298 24690
rect 4584 24774 9920 24784
rect 10500 24784 10510 28166
rect 10784 25716 10796 28256
rect 11020 25716 11032 28256
rect 12180 28256 12428 28718
rect 10784 25704 11032 25716
rect 11306 28166 11906 28176
rect 11306 24784 11316 28166
rect 10500 24774 11316 24784
rect 11896 24784 11906 28166
rect 12180 25716 12192 28256
rect 12416 25716 12428 28256
rect 13576 28256 13824 28718
rect 12180 25704 12428 25716
rect 12702 28166 13302 28176
rect 12702 24784 12712 28166
rect 11896 24774 12712 24784
rect 13292 24784 13302 28166
rect 13576 25716 13588 28256
rect 13812 25716 13824 28256
rect 14972 28256 15220 28718
rect 13576 25704 13824 25716
rect 14098 28166 14698 28176
rect 14098 24784 14108 28166
rect 13292 24774 14108 24784
rect 14688 24784 14698 28166
rect 14972 25716 14984 28256
rect 15208 25716 15220 28256
rect 16368 28256 16616 28718
rect 14972 25704 15220 25716
rect 15494 28166 16094 28176
rect 15494 24784 15504 28166
rect 14688 24774 15504 24784
rect 16084 24784 16094 28166
rect 16368 25716 16380 28256
rect 16604 25716 16616 28256
rect 17764 28256 18012 28718
rect 16368 25704 16616 25716
rect 16890 28166 17490 28176
rect 16890 24784 16900 28166
rect 16084 24774 16900 24784
rect 17480 24784 17490 28166
rect 17764 25716 17776 28256
rect 18000 25716 18012 28256
rect 19160 28256 19408 28718
rect 17764 25704 18012 25716
rect 18286 28166 18886 28176
rect 18286 24784 18296 28166
rect 17480 24774 18296 24784
rect 18876 24784 18886 28166
rect 19160 25716 19172 28256
rect 19396 25716 19408 28256
rect 20556 28256 20804 28718
rect 19160 25704 19408 25716
rect 19682 28166 20282 28176
rect 19682 24784 19692 28166
rect 18876 24774 19692 24784
rect 20272 24784 20282 28166
rect 20556 25716 20568 28256
rect 20792 25716 20804 28256
rect 21952 28256 22200 28718
rect 20556 25704 20804 25716
rect 21078 28166 21678 28176
rect 21078 24784 21088 28166
rect 20272 24774 21088 24784
rect 21668 24784 21678 28166
rect 21952 25716 21964 28256
rect 22188 25716 22200 28256
rect 23348 28256 23596 28718
rect 21952 25704 22200 25716
rect 22474 28166 23074 28176
rect 22474 24784 22484 28166
rect 21668 24774 22484 24784
rect 23064 24784 23074 28166
rect 23348 25716 23360 28256
rect 23584 25716 23596 28256
rect 24744 28256 24992 28718
rect 23348 25704 23596 25716
rect 23870 28166 24470 28176
rect 23870 24784 23880 28166
rect 23064 24774 23880 24784
rect 24460 24784 24470 28166
rect 24744 25716 24756 28256
rect 24980 25716 24992 28256
rect 26140 28256 26388 28718
rect 24744 25704 24992 25716
rect 25266 28166 25866 28176
rect 25266 24784 25276 28166
rect 24460 24774 25276 24784
rect 25856 24784 25866 28166
rect 26140 25716 26152 28256
rect 26376 25716 26388 28256
rect 27536 28256 27784 28718
rect 26140 25704 26388 25716
rect 26662 28166 27262 28176
rect 26662 24784 26672 28166
rect 25856 24774 26672 24784
rect 27252 24784 27262 28166
rect 27536 25716 27548 28256
rect 27772 25716 27784 28256
rect 28932 28256 29180 28718
rect 27536 25704 27784 25716
rect 28058 28166 28658 28176
rect 28058 24784 28068 28166
rect 27252 24774 28068 24784
rect 28648 24784 28658 28166
rect 28932 25716 28944 28256
rect 29168 25716 29180 28256
rect 30328 28256 30576 28718
rect 28932 25704 29180 25716
rect 29454 28166 30054 28176
rect 29454 24784 29464 28166
rect 28648 24774 29464 24784
rect 30044 24784 30054 28166
rect 30328 25716 30340 28256
rect 30564 25716 30576 28256
rect 31724 28256 31972 28718
rect 30328 25704 30576 25716
rect 30850 28166 31450 28176
rect 30850 24784 30860 28166
rect 30044 24774 30860 24784
rect 31440 24784 31450 28166
rect 31724 25716 31736 28256
rect 31960 25716 31972 28256
rect 33120 28256 33368 28718
rect 31724 25704 31972 25716
rect 32246 28166 32846 28176
rect 32246 24784 32256 28166
rect 31440 24774 32256 24784
rect 32836 24784 32846 28166
rect 33120 25716 33132 28256
rect 33356 25716 33368 28256
rect 34516 28256 34764 28718
rect 33120 25704 33368 25716
rect 33642 28166 34242 28176
rect 33642 24784 33652 28166
rect 32836 24774 33652 24784
rect 34232 24784 34242 28166
rect 34516 25716 34528 28256
rect 34752 25716 34764 28256
rect 35912 28256 36160 28718
rect 34516 25704 34764 25716
rect 35038 28166 35638 28176
rect 35038 24784 35048 28166
rect 34232 24774 35048 24784
rect 35628 24784 35638 28166
rect 35912 25716 35924 28256
rect 36148 25716 36160 28256
rect 37308 28256 37556 28718
rect 35912 25704 36160 25716
rect 36434 28166 37034 28176
rect 36434 24784 36444 28166
rect 35628 24774 36444 24784
rect 37024 24784 37034 28166
rect 37308 25716 37320 28256
rect 37544 25716 37556 28256
rect 38704 28256 38952 28718
rect 37308 25704 37556 25716
rect 37830 28166 38430 28176
rect 37830 24784 37840 28166
rect 37024 24774 37840 24784
rect 38420 24784 38430 28166
rect 38704 25716 38716 28256
rect 38940 25716 38952 28256
rect 40100 28256 40348 28718
rect 38704 25704 38952 25716
rect 39226 28166 39826 28176
rect 39226 24784 39236 28166
rect 38420 24774 39236 24784
rect 39816 24784 39826 28166
rect 40100 25716 40112 28256
rect 40336 25716 40348 28256
rect 41496 28256 41744 28718
rect 40100 25704 40348 25716
rect 40622 28166 41222 28176
rect 40622 24784 40632 28166
rect 39816 24774 40632 24784
rect 41212 24784 41222 28166
rect 41496 25716 41508 28256
rect 41732 25716 41744 28256
rect 42892 28256 43140 28718
rect 41496 25704 41744 25716
rect 42018 28166 42618 28176
rect 42018 24784 42028 28166
rect 41212 24774 42028 24784
rect 42608 24784 42618 28166
rect 42892 25716 42904 28256
rect 43128 25716 43140 28256
rect 44288 28256 44536 28718
rect 42892 25704 43140 25716
rect 43414 28166 44014 28176
rect 43414 24784 43424 28166
rect 42608 24774 43424 24784
rect 44004 24784 44014 28166
rect 44288 25716 44300 28256
rect 44524 25716 44536 28256
rect 45684 28256 45932 28718
rect 44288 25704 44536 25716
rect 44810 28166 45410 28176
rect 44810 24784 44820 28166
rect 44004 24774 44820 24784
rect 45400 24784 45410 28166
rect 45684 25716 45696 28256
rect 45920 25716 45932 28256
rect 47080 28256 47328 28718
rect 45684 25704 45932 25716
rect 46206 28166 46806 28176
rect 46206 24784 46216 28166
rect 45400 24774 46216 24784
rect 46796 24784 46806 28166
rect 47080 25716 47092 28256
rect 47316 25716 47328 28256
rect 48476 28256 48724 28718
rect 47080 25704 47328 25716
rect 47602 28166 48202 28176
rect 47602 24784 47612 28166
rect 46796 24774 47612 24784
rect 48192 24784 48202 28166
rect 48476 25716 48488 28256
rect 48712 25716 48724 28256
rect 49872 28256 50120 28718
rect 48476 25704 48724 25716
rect 48998 28166 49598 28176
rect 48998 24784 49008 28166
rect 48192 24774 49008 24784
rect 49588 24784 49598 28166
rect 49872 25716 49884 28256
rect 50108 25716 50120 28256
rect 49872 25704 50120 25716
rect 50394 28166 50994 28176
rect 50394 24784 50404 28166
rect 49588 24774 50404 24784
rect 50984 24784 50994 28166
rect 50984 24774 70094 24784
rect -1134 24446 -534 24448
rect 262 24446 862 24448
rect 1658 24446 2258 24448
rect 3054 24446 3654 24448
rect -2992 24438 3654 24446
rect -2992 23856 -1228 24438
rect 3618 23856 3654 24438
rect 4584 24394 4642 24774
rect 70084 24394 70094 24774
rect 4584 24384 70094 24394
rect 4624 24284 4688 24384
rect 4940 24284 5004 24384
rect 5256 24284 5320 24384
rect 5572 24284 5636 24384
rect 5888 24284 5952 24384
rect 6204 24284 6268 24384
rect 6520 24284 6584 24384
rect 6836 24284 6900 24384
rect 7152 24284 7216 24384
rect 7468 24284 7532 24384
rect 7784 24284 7848 24384
rect 8100 24284 8164 24384
rect 8416 24284 8480 24384
rect 8732 24284 8796 24384
rect 9048 24284 9112 24384
rect 9364 24284 9428 24384
rect 9680 24284 9744 24384
rect 9996 24284 10060 24384
rect 10312 24284 10376 24384
rect 10628 24284 10692 24384
rect 10944 24284 11008 24384
rect 11260 24284 11324 24384
rect 11576 24284 11640 24384
rect 11892 24284 11956 24384
rect 12208 24284 12272 24384
rect 12524 24284 12588 24384
rect 12840 24284 12904 24384
rect 13156 24284 13220 24384
rect 13472 24284 13536 24384
rect 13788 24284 13852 24384
rect 14104 24284 14168 24384
rect 14420 24284 14484 24384
rect 14736 24284 14800 24384
rect 15052 24284 15116 24384
rect 15368 24284 15432 24384
rect 15684 24284 15748 24384
rect 16000 24284 16064 24384
rect 16316 24284 16380 24384
rect 16632 24284 16696 24384
rect 16948 24284 17012 24384
rect 17264 24284 17328 24384
rect 17778 24284 17842 24384
rect 18094 24284 18158 24384
rect 18410 24284 18474 24384
rect 18726 24284 18790 24384
rect 19042 24284 19106 24384
rect 19358 24284 19422 24384
rect 19674 24284 19738 24384
rect 19990 24284 20054 24384
rect 20306 24284 20370 24384
rect 20622 24284 20686 24384
rect 20938 24284 21002 24384
rect 21254 24284 21318 24384
rect 21570 24284 21634 24384
rect 21886 24284 21950 24384
rect 22202 24284 22266 24384
rect 22518 24284 22582 24384
rect 22834 24284 22898 24384
rect 23150 24284 23214 24384
rect 23466 24284 23530 24384
rect 23782 24284 23846 24384
rect 24098 24284 24162 24384
rect 24414 24284 24478 24384
rect 24730 24284 24794 24384
rect 25046 24284 25110 24384
rect 25362 24284 25426 24384
rect 25678 24284 25742 24384
rect 25994 24284 26058 24384
rect 26310 24284 26374 24384
rect 26626 24284 26690 24384
rect 26942 24284 27006 24384
rect 27258 24284 27322 24384
rect 27574 24284 27638 24384
rect 27890 24284 27954 24384
rect 28206 24284 28270 24384
rect 28522 24284 28586 24384
rect 28838 24284 28902 24384
rect 29154 24284 29218 24384
rect 29470 24284 29534 24384
rect 29786 24284 29850 24384
rect 30102 24284 30166 24384
rect 30418 24284 30482 24384
rect 30932 24284 30996 24384
rect 31248 24284 31312 24384
rect 31564 24284 31628 24384
rect 31880 24284 31944 24384
rect 32196 24284 32260 24384
rect 32512 24284 32576 24384
rect 32828 24284 32892 24384
rect 33144 24284 33208 24384
rect 33460 24284 33524 24384
rect 33776 24284 33840 24384
rect 34092 24284 34156 24384
rect 34408 24284 34472 24384
rect 34724 24284 34788 24384
rect 35040 24284 35104 24384
rect 35356 24284 35420 24384
rect 35672 24284 35736 24384
rect 35988 24284 36052 24384
rect 36304 24284 36368 24384
rect 36620 24284 36684 24384
rect 36936 24284 37000 24384
rect 37252 24284 37316 24384
rect 37568 24284 37632 24384
rect 37884 24284 37948 24384
rect 38200 24284 38264 24384
rect 38516 24284 38580 24384
rect 38832 24284 38896 24384
rect 39148 24284 39212 24384
rect 39464 24284 39528 24384
rect 39780 24284 39844 24384
rect 40096 24284 40160 24384
rect 40412 24284 40476 24384
rect 40728 24284 40792 24384
rect 41044 24284 41108 24384
rect 41360 24284 41424 24384
rect 41676 24284 41740 24384
rect 41992 24284 42056 24384
rect 42308 24284 42372 24384
rect 42624 24284 42688 24384
rect 42940 24284 43004 24384
rect 43256 24284 43320 24384
rect 43572 24284 43636 24384
rect 44086 24284 44150 24384
rect 44402 24284 44466 24384
rect 44718 24284 44782 24384
rect 45034 24284 45098 24384
rect 45350 24284 45414 24384
rect 45666 24284 45730 24384
rect 45982 24284 46046 24384
rect 46298 24284 46362 24384
rect 46614 24284 46678 24384
rect 46930 24284 46994 24384
rect 47246 24284 47310 24384
rect 47562 24284 47626 24384
rect 47878 24284 47942 24384
rect 48194 24284 48258 24384
rect 48510 24284 48574 24384
rect 48826 24284 48890 24384
rect 49142 24284 49206 24384
rect 49458 24284 49522 24384
rect 49774 24284 49838 24384
rect 50090 24284 50154 24384
rect 50406 24284 50470 24384
rect 50722 24284 50786 24384
rect 51038 24284 51102 24384
rect 51354 24284 51418 24384
rect 51670 24284 51734 24384
rect 51986 24284 52050 24384
rect 52302 24284 52366 24384
rect 52618 24284 52682 24384
rect 52934 24284 52998 24384
rect 53250 24284 53314 24384
rect 53566 24284 53630 24384
rect 53882 24284 53946 24384
rect 54198 24284 54262 24384
rect 54514 24284 54578 24384
rect 54830 24284 54894 24384
rect 55146 24284 55210 24384
rect 55462 24284 55526 24384
rect 55778 24284 55842 24384
rect 56094 24284 56158 24384
rect 56410 24284 56474 24384
rect 56726 24284 56790 24384
rect 57240 24284 57304 24384
rect 57556 24284 57620 24384
rect 57872 24284 57936 24384
rect 58188 24284 58252 24384
rect 58504 24284 58568 24384
rect 58820 24284 58884 24384
rect 59136 24284 59200 24384
rect 59452 24284 59516 24384
rect 59768 24284 59832 24384
rect 60084 24284 60148 24384
rect 60400 24284 60464 24384
rect 60716 24284 60780 24384
rect 61032 24284 61096 24384
rect 61348 24284 61412 24384
rect 61664 24284 61728 24384
rect 61980 24284 62044 24384
rect 62296 24284 62360 24384
rect 62612 24284 62676 24384
rect 62928 24284 62992 24384
rect 63244 24284 63308 24384
rect 63560 24284 63624 24384
rect 63876 24284 63940 24384
rect 64192 24284 64256 24384
rect 64508 24284 64572 24384
rect 64824 24284 64888 24384
rect 65140 24284 65204 24384
rect 65456 24284 65520 24384
rect 65772 24284 65836 24384
rect 66088 24284 66152 24384
rect 66404 24284 66468 24384
rect 66720 24284 66784 24384
rect 67036 24284 67100 24384
rect 67352 24284 67416 24384
rect 67668 24284 67732 24384
rect 67984 24284 68048 24384
rect 68300 24284 68364 24384
rect 68616 24284 68680 24384
rect 68932 24284 68996 24384
rect 69248 24284 69312 24384
rect 69564 24284 69628 24384
rect 69880 24284 69944 24384
rect -2992 23846 3654 23856
rect 3165 23331 4181 23381
rect 3165 22941 3703 23331
rect 4093 22941 4181 23331
rect 3165 22791 4181 22941
rect 3165 19059 3755 22791
rect -3007 19035 3755 19059
rect -3007 18645 -2963 19035
rect -2573 18645 3755 19035
rect -3007 18469 3755 18645
rect 1305 15597 1895 18469
rect -17826 4066 -13826 12596
rect -3880 11686 -3870 12886
rect -3290 11686 -3280 12886
rect -3880 11676 -3280 11686
rect -1457 15007 1895 15597
rect -1457 8071 -867 15007
rect 4782 14276 4846 14372
rect 5098 14276 5162 14372
rect 5414 14276 5478 14372
rect 5730 14276 5794 14372
rect 6046 14276 6110 14372
rect 6362 14276 6426 14372
rect 6678 14276 6742 14372
rect 6994 14276 7058 14372
rect 7310 14276 7374 14372
rect 7626 14276 7690 14372
rect 7942 14276 8006 14372
rect 8258 14276 8322 14372
rect 8574 14276 8638 14372
rect 8890 14276 8954 14372
rect 9206 14276 9270 14372
rect 9522 14276 9586 14372
rect 9838 14276 9902 14372
rect 10154 14276 10218 14372
rect 10470 14276 10534 14372
rect 10786 14276 10850 14372
rect 11102 14276 11166 14372
rect 11418 14276 11482 14372
rect 11734 14276 11798 14372
rect 12050 14276 12114 14372
rect 12366 14276 12430 14372
rect 12682 14276 12746 14372
rect 12998 14276 13062 14372
rect 13314 14276 13378 14372
rect 13630 14276 13694 14372
rect 13946 14276 14010 14372
rect 14262 14276 14326 14372
rect 14578 14276 14642 14372
rect 14894 14276 14958 14372
rect 15210 14276 15274 14372
rect 15526 14276 15590 14372
rect 15842 14276 15906 14372
rect 16158 14276 16222 14372
rect 16474 14276 16538 14372
rect 16790 14276 16854 14372
rect 17106 14276 17170 14372
rect 17936 14276 18000 14372
rect 18252 14276 18316 14372
rect 18568 14276 18632 14372
rect 18884 14276 18948 14372
rect 19200 14276 19264 14372
rect 19516 14276 19580 14372
rect 19832 14276 19896 14372
rect 20148 14276 20212 14372
rect 20464 14276 20528 14372
rect 20780 14276 20844 14372
rect 21096 14276 21160 14372
rect 21412 14276 21476 14372
rect 21728 14276 21792 14372
rect 22044 14276 22108 14372
rect 22360 14276 22424 14372
rect 22676 14276 22740 14372
rect 22992 14276 23056 14372
rect 23308 14276 23372 14372
rect 23624 14276 23688 14372
rect 23940 14276 24004 14372
rect 24256 14276 24320 14372
rect 24572 14276 24636 14372
rect 24888 14276 24952 14372
rect 25204 14276 25268 14372
rect 25520 14276 25584 14372
rect 25836 14276 25900 14372
rect 26152 14276 26216 14372
rect 26468 14276 26532 14372
rect 26784 14276 26848 14372
rect 27100 14276 27164 14372
rect 27416 14276 27480 14372
rect 27732 14276 27796 14372
rect 28048 14276 28112 14372
rect 28364 14276 28428 14372
rect 28680 14276 28744 14372
rect 28996 14276 29060 14372
rect 29312 14276 29376 14372
rect 29628 14276 29692 14372
rect 29944 14276 30008 14372
rect 30260 14276 30324 14372
rect 31090 14276 31154 14372
rect 31406 14276 31470 14372
rect 31722 14276 31786 14372
rect 32038 14276 32102 14372
rect 32354 14276 32418 14372
rect 32670 14276 32734 14372
rect 32986 14276 33050 14372
rect 33302 14276 33366 14372
rect 33618 14276 33682 14372
rect 33934 14276 33998 14372
rect 34250 14276 34314 14372
rect 34566 14276 34630 14372
rect 34882 14276 34946 14372
rect 35198 14276 35262 14372
rect 35514 14276 35578 14372
rect 35830 14276 35894 14372
rect 36146 14276 36210 14372
rect 36462 14276 36526 14372
rect 36778 14276 36842 14372
rect 37094 14276 37158 14372
rect 37410 14276 37474 14372
rect 37726 14276 37790 14372
rect 38042 14276 38106 14372
rect 38358 14276 38422 14372
rect 38674 14276 38738 14372
rect 38990 14276 39054 14372
rect 39306 14276 39370 14372
rect 39622 14276 39686 14372
rect 39938 14276 40002 14372
rect 40254 14276 40318 14372
rect 40570 14276 40634 14372
rect 40886 14276 40950 14372
rect 41202 14276 41266 14372
rect 41518 14276 41582 14372
rect 41834 14276 41898 14372
rect 42150 14276 42214 14372
rect 42466 14276 42530 14372
rect 42782 14276 42846 14372
rect 43098 14276 43162 14372
rect 43414 14276 43478 14372
rect 44244 14276 44308 14372
rect 44560 14276 44624 14372
rect 44876 14276 44940 14372
rect 45192 14276 45256 14372
rect 45508 14276 45572 14372
rect 45824 14276 45888 14372
rect 46140 14276 46204 14372
rect 46456 14276 46520 14372
rect 46772 14276 46836 14372
rect 47088 14276 47152 14372
rect 47404 14276 47468 14372
rect 47720 14276 47784 14372
rect 48036 14276 48100 14372
rect 48352 14276 48416 14372
rect 48668 14276 48732 14372
rect 48984 14276 49048 14372
rect 49300 14276 49364 14372
rect 49616 14276 49680 14372
rect 49932 14276 49996 14372
rect 50248 14276 50312 14372
rect 50564 14276 50628 14372
rect 50880 14276 50944 14372
rect 51196 14276 51260 14372
rect 51512 14276 51576 14372
rect 51828 14276 51892 14372
rect 52144 14276 52208 14372
rect 52460 14276 52524 14372
rect 52776 14276 52840 14372
rect 53092 14276 53156 14372
rect 53408 14276 53472 14372
rect 53724 14276 53788 14372
rect 54040 14276 54104 14372
rect 54356 14276 54420 14372
rect 54672 14276 54736 14372
rect 54988 14276 55052 14372
rect 55304 14276 55368 14372
rect 55620 14276 55684 14372
rect 55936 14276 56000 14372
rect 56252 14276 56316 14372
rect 56568 14276 56632 14372
rect 57398 14276 57462 14372
rect 57714 14276 57778 14372
rect 58030 14276 58094 14372
rect 58346 14276 58410 14372
rect 58662 14276 58726 14372
rect 58978 14276 59042 14372
rect 59294 14276 59358 14372
rect 59610 14276 59674 14372
rect 59926 14276 59990 14372
rect 60242 14276 60306 14372
rect 60558 14276 60622 14372
rect 60874 14276 60938 14372
rect 61190 14276 61254 14372
rect 61506 14276 61570 14372
rect 61822 14276 61886 14372
rect 62138 14276 62202 14372
rect 62454 14276 62518 14372
rect 62770 14276 62834 14372
rect 63086 14276 63150 14372
rect 63402 14276 63466 14372
rect 63718 14276 63782 14372
rect 64034 14276 64098 14372
rect 64350 14276 64414 14372
rect 64666 14276 64730 14372
rect 64982 14276 65046 14372
rect 65298 14276 65362 14372
rect 65614 14276 65678 14372
rect 65930 14276 65994 14372
rect 66246 14276 66310 14372
rect 66562 14276 66626 14372
rect 66878 14276 66942 14372
rect 67194 14276 67258 14372
rect 67510 14276 67574 14372
rect 67826 14276 67890 14372
rect 68142 14276 68206 14372
rect 68458 14276 68522 14372
rect 68774 14276 68838 14372
rect 69090 14276 69154 14372
rect 69406 14276 69470 14372
rect 69722 14276 69786 14372
rect 4568 14182 69954 14276
rect 4568 12856 4662 14182
rect 69856 12856 69954 14182
rect 4568 12744 69954 12856
rect -1457 7481 1928 8071
rect 1338 4844 1928 7481
rect 1338 4440 1938 4844
rect 1146 4430 3386 4440
rect 1146 4420 1370 4430
rect 1146 4066 1362 4420
rect -17826 66 1362 4066
rect 3376 124 3386 4430
rect 3376 66 3406 124
rect 1336 22 3406 66
<< via3 >>
rect -17422 29110 -16842 29690
rect -16222 29110 -15642 29690
rect -15022 29110 -14442 29690
rect -13822 29110 -13242 29690
rect -12622 29110 -12042 29690
rect -11422 29110 -10842 29690
rect -10222 29110 -9642 29690
rect -9022 29110 -8442 29690
rect -7822 29110 -7242 29690
rect -6622 29110 -6042 29690
rect -5422 29110 -4842 29690
rect -3870 28490 -3290 29690
rect 4642 24394 70084 24774
rect -3870 11686 -3290 12886
rect 4662 12856 69856 14182
rect 1370 4420 3376 4430
rect 1362 4048 1370 4420
rect 1370 4048 3362 4420
rect 1362 3740 1376 4048
rect 1376 3740 3362 4048
rect 3362 3740 3376 4420
rect 1362 66 3376 3740
<< metal4 >>
rect -17432 29690 -3280 29700
rect -17432 29110 -17422 29690
rect -16842 29110 -16222 29690
rect -15642 29110 -15022 29690
rect -14442 29110 -13822 29690
rect -13242 29110 -12622 29690
rect -12042 29110 -11422 29690
rect -10842 29110 -10222 29690
rect -9642 29110 -9022 29690
rect -8442 29110 -7822 29690
rect -7242 29110 -6622 29690
rect -6042 29110 -5422 29690
rect -4842 29110 -3870 29690
rect -17432 29100 -3870 29110
rect -3880 28490 -3870 29100
rect -3290 28490 -3280 29690
rect -3880 12886 -3280 28490
rect 4584 24872 70094 24920
rect 4584 24428 4636 24872
rect 70042 24774 70094 24872
rect 4584 24394 4642 24428
rect 70084 24394 70094 24774
rect 4584 24384 70094 24394
rect -3880 11686 -3870 12886
rect -3290 11686 -3280 12886
rect 4568 14182 69954 14276
rect 4568 12856 4662 14182
rect 69856 12856 69954 14182
rect 4568 12744 69954 12856
rect -3880 11676 -3280 11686
rect 1336 4430 3386 4440
rect 1336 4420 1370 4430
rect 1336 66 1362 4420
rect 3376 124 3386 4430
rect 3376 66 3406 124
rect 1336 22 3406 66
<< via4 >>
rect 4636 24774 70042 24872
rect 4636 24428 4642 24774
rect 4642 24428 70042 24774
rect 4662 12856 69856 14182
rect 1362 66 3362 4420
<< metal5 >>
rect 4584 24872 70094 24920
rect 4584 24428 4636 24872
rect 70042 24428 70094 24872
rect 4584 24384 70094 24428
rect 4568 14182 69954 14276
rect 4568 12856 4662 14182
rect 69856 12856 69954 14182
rect 4568 11212 69954 12856
rect 1338 4440 3408 4480
rect 1336 4420 3408 4440
rect 1336 66 1362 4420
rect 3362 4374 3408 4420
rect 4568 4374 7632 11212
rect 3362 1310 7632 4374
rect 3362 66 3408 1310
rect 1336 22 3406 66
use large_nmos_g5d10  large_nmos_g5d10_0
timestamp 1664842101
transform 1 0 30830 0 1 19394
box -124 -66 13030 4890
use large_nmos_g5d10  large_nmos_g5d10_1
timestamp 1664842101
transform 1 0 43984 0 1 19394
box -124 -66 13030 4890
use large_nmos_g5d10  large_nmos_g5d10_2
timestamp 1664842101
transform 1 0 57138 0 1 19394
box -124 -66 13030 4890
use large_nmos_g5d10  large_nmos_g5d10_3
timestamp 1664842101
transform 1 0 4522 0 1 14438
box -124 -66 13030 4890
use large_nmos_g5d10  large_nmos_g5d10_4
timestamp 1664842101
transform 1 0 4522 0 1 19394
box -124 -66 13030 4890
use large_nmos_g5d10  large_nmos_g5d10_5
timestamp 1664842101
transform 1 0 17676 0 1 19394
box -124 -66 13030 4890
use large_nmos_g5d10  large_nmos_g5d10_6
timestamp 1664842101
transform 1 0 17676 0 1 14438
box -124 -66 13030 4890
use large_nmos_g5d10  large_nmos_g5d10_7
timestamp 1664842101
transform 1 0 30830 0 1 14438
box -124 -66 13030 4890
use large_nmos_g5d10  large_nmos_g5d10_8
timestamp 1664842101
transform 1 0 43984 0 1 14438
box -124 -66 13030 4890
use large_nmos_g5d10  large_nmos_g5d10_9
timestamp 1664842101
transform 1 0 57138 0 1 14438
box -124 -66 13030 4890
use sky130_fd_pr__diode_pd2nw_11v0_6YHF4V  sky130_fd_pr__diode_pd2nw_11v0_6YHF4V_0
timestamp 1665170787
transform 1 0 1260 0 1 27596
box -2972 -2972 2972 2972
use sky130_fd_pr__diode_pd2nw_11v0_VFE9GT  sky130_fd_pr__diode_pd2nw_11v0_VFE9GT_0
timestamp 1667507583
transform 1 0 30452 0 1 27034
box -21120 -1576 21120 1576
use sky130_fd_pr__nfet_g5v0d10v5_U5GC69  sky130_fd_pr__nfet_g5v0d10v5_U5GC69_0
timestamp 1664842101
transform 1 0 1995 0 1 11707
box -1779 -1753 1779 1753
use sky130_fd_pr__rf_npn_05v5_W1p00L2p00  sky130_fd_pr__rf_npn_05v5_W1p00L2p00_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1661821916
transform 1 0 -4940 0 1 8112
box 0 0 1724 1924
use sky130_fd_pr__rf_npn_05v5_W1p00L2p00  sky130_fd_pr__rf_npn_05v5_W1p00L2p00_1
array 0 3 1406 0 3 1606
timestamp 1661821916
transform 1 0 -12922 0 1 5364
box 0 0 1724 1924
use sky130_fd_pr__rf_npn_05v5_W1p00L2p00  sky130_fd_pr__rf_npn_05v5_W1p00L2p00_2
array 0 9 1406 0 9 1606
timestamp 1661821916
transform 1 0 -18550 0 1 13256
box 0 0 1724 1924
<< labels >>
rlabel metal3 s 6794 24746 6794 24746 1 VsMOS
rlabel metal1 3928 14760 3928 14760 1 VpMOS
rlabel metal1 s -17890 29920 -17890 29920 1 VsBJT
rlabel metal1 -6444 8138 -6444 8138 1 VpBJT
rlabel metal5 6440 3684 6440 3684 1 Ground
rlabel via2 10146 28742 10146 28742 1 Vo
<< end >>
