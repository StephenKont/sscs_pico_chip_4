magic
tech sky130A
timestamp 1669944869
<< pwell >>
rect -1172 -1129 1172 1129
<< mvnmos >>
rect -1058 -1000 -658 1000
rect -629 -1000 -229 1000
rect -200 -1000 200 1000
rect 229 -1000 629 1000
rect 658 -1000 1058 1000
<< mvndiff >>
rect -1087 994 -1058 1000
rect -1087 -994 -1081 994
rect -1064 -994 -1058 994
rect -1087 -1000 -1058 -994
rect -658 994 -629 1000
rect -658 -994 -652 994
rect -635 -994 -629 994
rect -658 -1000 -629 -994
rect -229 994 -200 1000
rect -229 -994 -223 994
rect -206 -994 -200 994
rect -229 -1000 -200 -994
rect 200 994 229 1000
rect 200 -994 206 994
rect 223 -994 229 994
rect 200 -1000 229 -994
rect 629 994 658 1000
rect 629 -994 635 994
rect 652 -994 658 994
rect 629 -1000 658 -994
rect 1058 994 1087 1000
rect 1058 -994 1064 994
rect 1081 -994 1087 994
rect 1058 -1000 1087 -994
<< mvndiffc >>
rect -1081 -994 -1064 994
rect -652 -994 -635 994
rect -223 -994 -206 994
rect 206 -994 223 994
rect 635 -994 652 994
rect 1064 -994 1081 994
<< mvpsubdiff >>
rect -1154 1105 1154 1111
rect -1154 1088 -1100 1105
rect 1100 1088 1154 1105
rect -1154 1082 1154 1088
rect -1154 1057 -1125 1082
rect -1154 -1057 -1148 1057
rect -1131 -1057 -1125 1057
rect 1125 1057 1154 1082
rect -1154 -1082 -1125 -1057
rect 1125 -1057 1131 1057
rect 1148 -1057 1154 1057
rect 1125 -1082 1154 -1057
rect -1154 -1088 1154 -1082
rect -1154 -1105 -1100 -1088
rect 1100 -1105 1154 -1088
rect -1154 -1111 1154 -1105
<< mvpsubdiffcont >>
rect -1100 1088 1100 1105
rect -1148 -1057 -1131 1057
rect 1131 -1057 1148 1057
rect -1100 -1105 1100 -1088
<< poly >>
rect -1058 1036 -658 1044
rect -1058 1019 -1050 1036
rect -666 1019 -658 1036
rect -1058 1000 -658 1019
rect -629 1036 -229 1044
rect -629 1019 -621 1036
rect -237 1019 -229 1036
rect -629 1000 -229 1019
rect -200 1036 200 1044
rect -200 1019 -192 1036
rect 192 1019 200 1036
rect -200 1000 200 1019
rect 229 1036 629 1044
rect 229 1019 237 1036
rect 621 1019 629 1036
rect 229 1000 629 1019
rect 658 1036 1058 1044
rect 658 1019 666 1036
rect 1050 1019 1058 1036
rect 658 1000 1058 1019
rect -1058 -1019 -658 -1000
rect -1058 -1036 -1050 -1019
rect -666 -1036 -658 -1019
rect -1058 -1044 -658 -1036
rect -629 -1019 -229 -1000
rect -629 -1036 -621 -1019
rect -237 -1036 -229 -1019
rect -629 -1044 -229 -1036
rect -200 -1019 200 -1000
rect -200 -1036 -192 -1019
rect 192 -1036 200 -1019
rect -200 -1044 200 -1036
rect 229 -1019 629 -1000
rect 229 -1036 237 -1019
rect 621 -1036 629 -1019
rect 229 -1044 629 -1036
rect 658 -1019 1058 -1000
rect 658 -1036 666 -1019
rect 1050 -1036 1058 -1019
rect 658 -1044 1058 -1036
<< polycont >>
rect -1050 1019 -666 1036
rect -621 1019 -237 1036
rect -192 1019 192 1036
rect 237 1019 621 1036
rect 666 1019 1050 1036
rect -1050 -1036 -666 -1019
rect -621 -1036 -237 -1019
rect -192 -1036 192 -1019
rect 237 -1036 621 -1019
rect 666 -1036 1050 -1019
<< locali >>
rect -1148 1088 -1100 1105
rect 1100 1088 1148 1105
rect -1148 1057 -1131 1088
rect 1131 1057 1148 1088
rect -1058 1019 -1050 1036
rect -666 1019 -658 1036
rect -629 1019 -621 1036
rect -237 1019 -229 1036
rect -200 1019 -192 1036
rect 192 1019 200 1036
rect 229 1019 237 1036
rect 621 1019 629 1036
rect 658 1019 666 1036
rect 1050 1019 1058 1036
rect -1081 994 -1064 1002
rect -1131 500 -1081 600
rect -1131 100 -1081 200
rect -1131 -300 -1081 -200
rect -1131 -700 -1081 -600
rect -652 994 -635 1002
rect -1064 500 -652 600
rect -1064 100 -652 200
rect -1064 -300 -652 -200
rect -1064 -700 -652 -600
rect -1081 -1002 -1064 -994
rect -223 994 -206 1002
rect -635 500 -223 600
rect -635 100 -223 200
rect -635 -300 -223 -200
rect -635 -700 -223 -600
rect -652 -1002 -635 -994
rect 206 994 223 1002
rect -206 500 206 600
rect -206 100 206 200
rect -206 -300 206 -200
rect -206 -700 206 -600
rect -223 -1002 -206 -994
rect 635 994 652 1002
rect 223 500 635 600
rect 223 100 635 200
rect 223 -300 635 -200
rect 223 -700 635 -600
rect 206 -1002 223 -994
rect 1064 994 1081 1002
rect 652 500 1064 600
rect 652 100 1064 200
rect 652 -300 1064 -200
rect 652 -700 1064 -600
rect 635 -1002 652 -994
rect 1081 500 1131 600
rect 1081 100 1131 200
rect 1081 -300 1131 -200
rect 1081 -700 1131 -600
rect 1064 -1002 1081 -994
rect -1058 -1036 -1050 -1019
rect -666 -1036 -658 -1019
rect -629 -1036 -621 -1019
rect -237 -1036 -229 -1019
rect -200 -1036 -192 -1019
rect 192 -1036 200 -1019
rect 229 -1036 237 -1019
rect 621 -1036 629 -1019
rect 658 -1036 666 -1019
rect 1050 -1036 1058 -1019
rect -1148 -1088 -1131 -1057
rect 1131 -1088 1148 -1057
rect -1148 -1105 -1100 -1088
rect 1100 -1105 1148 -1088
<< viali >>
rect -1050 1019 -666 1036
rect -621 1019 -237 1036
rect -192 1019 192 1036
rect 237 1019 621 1036
rect 666 1019 1050 1036
rect -1081 -994 -1064 994
rect -652 -994 -635 994
rect -223 -994 -206 994
rect 206 -994 223 994
rect 635 -994 652 994
rect 1064 -994 1081 994
rect -1050 -1036 -666 -1019
rect -621 -1036 -237 -1019
rect -192 -1036 192 -1019
rect 237 -1036 621 -1019
rect 666 -1036 1050 -1019
<< metal1 >>
rect -1058 1069 1058 1072
rect -1058 1019 -1055 1069
rect 1055 1019 1058 1069
rect -1058 1016 1058 1019
rect -1084 994 -1061 1000
rect -1084 -994 -1081 994
rect -1064 -994 -1061 994
rect -1084 -1000 -1061 -994
rect -655 994 -632 1000
rect -655 -994 -652 994
rect -635 -994 -632 994
rect -655 -1000 -632 -994
rect -226 994 -203 1000
rect -226 -994 -223 994
rect -206 -994 -203 994
rect -226 -1000 -203 -994
rect 203 994 226 1000
rect 203 -994 206 994
rect 223 -994 226 994
rect 203 -1000 226 -994
rect 632 994 655 1000
rect 632 -994 635 994
rect 652 -994 655 994
rect 632 -1000 655 -994
rect 1061 994 1084 1000
rect 1061 -994 1064 994
rect 1081 -994 1084 994
rect 1061 -1000 1084 -994
rect -1058 -1019 1058 -1016
rect -1058 -1069 -1055 -1019
rect 1055 -1069 1058 -1019
rect -1058 -1072 1058 -1069
<< via1 >>
rect -1055 1036 1055 1069
rect -1055 1019 -1050 1036
rect -1050 1019 -666 1036
rect -666 1019 -621 1036
rect -621 1019 -237 1036
rect -237 1019 -192 1036
rect -192 1019 192 1036
rect 192 1019 237 1036
rect 237 1019 621 1036
rect 621 1019 666 1036
rect 666 1019 1050 1036
rect 1050 1019 1055 1036
rect -1055 -1036 -1050 -1019
rect -1050 -1036 -666 -1019
rect -666 -1036 -621 -1019
rect -621 -1036 -237 -1019
rect -237 -1036 -192 -1019
rect -192 -1036 192 -1019
rect 192 -1036 237 -1019
rect 237 -1036 621 -1019
rect 621 -1036 666 -1019
rect 666 -1036 1050 -1019
rect 1050 -1036 1055 -1019
rect -1055 -1069 1055 -1036
<< metal2 >>
rect -1058 1069 1058 1072
rect -1058 1019 -1055 1069
rect 1055 1019 1058 1069
rect -1058 1016 1058 1019
rect -1058 -1019 1058 -1016
rect -1058 -1069 -1055 -1019
rect 1055 -1069 1058 -1019
rect -1058 -1072 1058 -1069
<< properties >>
string FIXED_BBOX -1139 -1096 1139 1096
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 20 l 4 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
