magic
tech sky130A
magscale 1 2
timestamp 1668293870
<< pwell >>
rect -783 -410 783 410
<< nmos >>
rect -587 -200 -337 200
rect -279 -200 -29 200
rect 29 -200 279 200
rect 337 -200 587 200
<< ndiff >>
rect -645 188 -587 200
rect -645 -188 -633 188
rect -599 -188 -587 188
rect -645 -200 -587 -188
rect -337 188 -279 200
rect -337 -188 -325 188
rect -291 -188 -279 188
rect -337 -200 -279 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 279 188 337 200
rect 279 -188 291 188
rect 325 -188 337 188
rect 279 -200 337 -188
rect 587 188 645 200
rect 587 -188 599 188
rect 633 -188 645 188
rect 587 -200 645 -188
<< ndiffc >>
rect -633 -188 -599 188
rect -325 -188 -291 188
rect -17 -188 17 188
rect 291 -188 325 188
rect 599 -188 633 188
<< psubdiff >>
rect -747 340 -651 374
rect 651 340 747 374
rect -747 278 -713 340
rect 713 278 747 340
rect -747 -340 -713 -278
rect 713 -340 747 -278
rect -747 -374 -651 -340
rect 651 -374 747 -340
<< psubdiffcont >>
rect -651 340 651 374
rect -747 -278 -713 278
rect 713 -278 747 278
rect -651 -374 651 -340
<< poly >>
rect -587 272 -337 288
rect -587 238 -571 272
rect -353 238 -337 272
rect -587 200 -337 238
rect -279 272 -29 288
rect -279 238 -263 272
rect -45 238 -29 272
rect -279 200 -29 238
rect 29 272 279 288
rect 29 238 45 272
rect 263 238 279 272
rect 29 200 279 238
rect 337 272 587 288
rect 337 238 353 272
rect 571 238 587 272
rect 337 200 587 238
rect -587 -238 -337 -200
rect -587 -272 -571 -238
rect -353 -272 -337 -238
rect -587 -288 -337 -272
rect -279 -238 -29 -200
rect -279 -272 -263 -238
rect -45 -272 -29 -238
rect -279 -288 -29 -272
rect 29 -238 279 -200
rect 29 -272 45 -238
rect 263 -272 279 -238
rect 29 -288 279 -272
rect 337 -238 587 -200
rect 337 -272 353 -238
rect 571 -272 587 -238
rect 337 -288 587 -272
<< polycont >>
rect -571 238 -353 272
rect -263 238 -45 272
rect 45 238 263 272
rect 353 238 571 272
rect -571 -272 -353 -238
rect -263 -272 -45 -238
rect 45 -272 263 -238
rect 353 -272 571 -238
<< locali >>
rect -747 340 -651 374
rect 651 340 747 374
rect -747 278 -713 340
rect 713 278 747 340
rect -587 238 -571 272
rect -353 238 -337 272
rect -279 238 -263 272
rect -45 238 -29 272
rect 29 238 45 272
rect 263 238 279 272
rect 337 238 353 272
rect 571 238 587 272
rect -633 188 -599 204
rect -633 -204 -599 -188
rect -325 188 -291 204
rect -325 -204 -291 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 291 188 325 204
rect 291 -204 325 -188
rect 599 188 633 204
rect 599 -204 633 -188
rect -587 -272 -571 -238
rect -353 -272 -337 -238
rect -279 -272 -263 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 263 -272 279 -238
rect 337 -272 353 -238
rect 571 -272 587 -238
rect -747 -340 -713 -278
rect 713 -340 747 -278
rect -747 -374 -651 -340
rect 651 -374 747 -340
<< viali >>
rect -571 238 -353 272
rect -263 238 -45 272
rect 45 238 263 272
rect 353 238 571 272
rect -633 -188 -599 188
rect -325 -188 -291 188
rect -17 -188 17 188
rect 291 -188 325 188
rect 599 -188 633 188
rect -571 -272 -353 -238
rect -263 -272 -45 -238
rect 45 -272 263 -238
rect 353 -272 571 -238
<< metal1 >>
rect -583 272 -341 278
rect -583 238 -571 272
rect -353 238 -341 272
rect -583 232 -341 238
rect -275 272 -33 278
rect -275 238 -263 272
rect -45 238 -33 272
rect -275 232 -33 238
rect 33 272 275 278
rect 33 238 45 272
rect 263 238 275 272
rect 33 232 275 238
rect 341 272 583 278
rect 341 238 353 272
rect 571 238 583 272
rect 341 232 583 238
rect -639 188 -593 200
rect -639 -188 -633 188
rect -599 -188 -593 188
rect -639 -200 -593 -188
rect -331 188 -285 200
rect -331 -188 -325 188
rect -291 -188 -285 188
rect -331 -200 -285 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 285 188 331 200
rect 285 -188 291 188
rect 325 -188 331 188
rect 285 -200 331 -188
rect 593 188 639 200
rect 593 -188 599 188
rect 633 -188 639 188
rect 593 -200 639 -188
rect -583 -238 -341 -232
rect -583 -272 -571 -238
rect -353 -272 -341 -238
rect -583 -278 -341 -272
rect -275 -238 -33 -232
rect -275 -272 -263 -238
rect -45 -272 -33 -238
rect -275 -278 -33 -272
rect 33 -238 275 -232
rect 33 -272 45 -238
rect 263 -272 275 -238
rect 33 -278 275 -272
rect 341 -238 583 -232
rect 341 -272 353 -238
rect 571 -272 583 -238
rect 341 -278 583 -272
<< properties >>
string FIXED_BBOX -730 -357 730 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
