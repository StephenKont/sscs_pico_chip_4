magic
tech sky130A
timestamp 1665174684
<< nwell >>
rect -5235 -1396 5235 1396
<< pwell >>
rect -5325 1396 5325 1486
rect -5325 -1396 -5235 1396
rect 5235 -1396 5325 1396
rect -5325 -1486 5325 -1396
<< mvpsubdiff >>
rect -5307 1462 5307 1468
rect -5307 1445 -5253 1462
rect 5253 1445 5307 1462
rect -5307 1439 5307 1445
rect -5307 1414 -5278 1439
rect -5307 -1414 -5301 1414
rect -5284 -1414 -5278 1414
rect 5278 1414 5307 1439
rect -5307 -1439 -5278 -1414
rect 5278 -1414 5284 1414
rect 5301 -1414 5307 1414
rect 5278 -1439 5307 -1414
rect -5307 -1445 5307 -1439
rect -5307 -1462 -5253 -1445
rect 5253 -1462 5307 -1445
rect -5307 -1468 5307 -1462
<< mvnsubdiff >>
rect -5202 1357 -4570 1363
rect -5202 1340 -5148 1357
rect -4624 1340 -4570 1357
rect -5202 1334 -4570 1340
rect -5202 1309 -5173 1334
rect -5202 785 -5196 1309
rect -5179 785 -5173 1309
rect -4599 1309 -4570 1334
rect -5202 760 -5173 785
rect -4599 785 -4593 1309
rect -4576 785 -4570 1309
rect -4599 760 -4570 785
rect -5202 754 -4570 760
rect -5202 737 -5148 754
rect -4624 737 -4570 754
rect -5202 731 -4570 737
rect -4504 1357 -3872 1363
rect -4504 1340 -4450 1357
rect -3926 1340 -3872 1357
rect -4504 1334 -3872 1340
rect -4504 1309 -4475 1334
rect -4504 785 -4498 1309
rect -4481 785 -4475 1309
rect -3901 1309 -3872 1334
rect -4504 760 -4475 785
rect -3901 785 -3895 1309
rect -3878 785 -3872 1309
rect -3901 760 -3872 785
rect -4504 754 -3872 760
rect -4504 737 -4450 754
rect -3926 737 -3872 754
rect -4504 731 -3872 737
rect -3806 1357 -3174 1363
rect -3806 1340 -3752 1357
rect -3228 1340 -3174 1357
rect -3806 1334 -3174 1340
rect -3806 1309 -3777 1334
rect -3806 785 -3800 1309
rect -3783 785 -3777 1309
rect -3203 1309 -3174 1334
rect -3806 760 -3777 785
rect -3203 785 -3197 1309
rect -3180 785 -3174 1309
rect -3203 760 -3174 785
rect -3806 754 -3174 760
rect -3806 737 -3752 754
rect -3228 737 -3174 754
rect -3806 731 -3174 737
rect -3108 1357 -2476 1363
rect -3108 1340 -3054 1357
rect -2530 1340 -2476 1357
rect -3108 1334 -2476 1340
rect -3108 1309 -3079 1334
rect -3108 785 -3102 1309
rect -3085 785 -3079 1309
rect -2505 1309 -2476 1334
rect -3108 760 -3079 785
rect -2505 785 -2499 1309
rect -2482 785 -2476 1309
rect -2505 760 -2476 785
rect -3108 754 -2476 760
rect -3108 737 -3054 754
rect -2530 737 -2476 754
rect -3108 731 -2476 737
rect -2410 1357 -1778 1363
rect -2410 1340 -2356 1357
rect -1832 1340 -1778 1357
rect -2410 1334 -1778 1340
rect -2410 1309 -2381 1334
rect -2410 785 -2404 1309
rect -2387 785 -2381 1309
rect -1807 1309 -1778 1334
rect -2410 760 -2381 785
rect -1807 785 -1801 1309
rect -1784 785 -1778 1309
rect -1807 760 -1778 785
rect -2410 754 -1778 760
rect -2410 737 -2356 754
rect -1832 737 -1778 754
rect -2410 731 -1778 737
rect -1712 1357 -1080 1363
rect -1712 1340 -1658 1357
rect -1134 1340 -1080 1357
rect -1712 1334 -1080 1340
rect -1712 1309 -1683 1334
rect -1712 785 -1706 1309
rect -1689 785 -1683 1309
rect -1109 1309 -1080 1334
rect -1712 760 -1683 785
rect -1109 785 -1103 1309
rect -1086 785 -1080 1309
rect -1109 760 -1080 785
rect -1712 754 -1080 760
rect -1712 737 -1658 754
rect -1134 737 -1080 754
rect -1712 731 -1080 737
rect -1014 1357 -382 1363
rect -1014 1340 -960 1357
rect -436 1340 -382 1357
rect -1014 1334 -382 1340
rect -1014 1309 -985 1334
rect -1014 785 -1008 1309
rect -991 785 -985 1309
rect -411 1309 -382 1334
rect -1014 760 -985 785
rect -411 785 -405 1309
rect -388 785 -382 1309
rect -411 760 -382 785
rect -1014 754 -382 760
rect -1014 737 -960 754
rect -436 737 -382 754
rect -1014 731 -382 737
rect -316 1357 316 1363
rect -316 1340 -262 1357
rect 262 1340 316 1357
rect -316 1334 316 1340
rect -316 1309 -287 1334
rect -316 785 -310 1309
rect -293 785 -287 1309
rect 287 1309 316 1334
rect -316 760 -287 785
rect 287 785 293 1309
rect 310 785 316 1309
rect 287 760 316 785
rect -316 754 316 760
rect -316 737 -262 754
rect 262 737 316 754
rect -316 731 316 737
rect 382 1357 1014 1363
rect 382 1340 436 1357
rect 960 1340 1014 1357
rect 382 1334 1014 1340
rect 382 1309 411 1334
rect 382 785 388 1309
rect 405 785 411 1309
rect 985 1309 1014 1334
rect 382 760 411 785
rect 985 785 991 1309
rect 1008 785 1014 1309
rect 985 760 1014 785
rect 382 754 1014 760
rect 382 737 436 754
rect 960 737 1014 754
rect 382 731 1014 737
rect 1080 1357 1712 1363
rect 1080 1340 1134 1357
rect 1658 1340 1712 1357
rect 1080 1334 1712 1340
rect 1080 1309 1109 1334
rect 1080 785 1086 1309
rect 1103 785 1109 1309
rect 1683 1309 1712 1334
rect 1080 760 1109 785
rect 1683 785 1689 1309
rect 1706 785 1712 1309
rect 1683 760 1712 785
rect 1080 754 1712 760
rect 1080 737 1134 754
rect 1658 737 1712 754
rect 1080 731 1712 737
rect 1778 1357 2410 1363
rect 1778 1340 1832 1357
rect 2356 1340 2410 1357
rect 1778 1334 2410 1340
rect 1778 1309 1807 1334
rect 1778 785 1784 1309
rect 1801 785 1807 1309
rect 2381 1309 2410 1334
rect 1778 760 1807 785
rect 2381 785 2387 1309
rect 2404 785 2410 1309
rect 2381 760 2410 785
rect 1778 754 2410 760
rect 1778 737 1832 754
rect 2356 737 2410 754
rect 1778 731 2410 737
rect 2476 1357 3108 1363
rect 2476 1340 2530 1357
rect 3054 1340 3108 1357
rect 2476 1334 3108 1340
rect 2476 1309 2505 1334
rect 2476 785 2482 1309
rect 2499 785 2505 1309
rect 3079 1309 3108 1334
rect 2476 760 2505 785
rect 3079 785 3085 1309
rect 3102 785 3108 1309
rect 3079 760 3108 785
rect 2476 754 3108 760
rect 2476 737 2530 754
rect 3054 737 3108 754
rect 2476 731 3108 737
rect 3174 1357 3806 1363
rect 3174 1340 3228 1357
rect 3752 1340 3806 1357
rect 3174 1334 3806 1340
rect 3174 1309 3203 1334
rect 3174 785 3180 1309
rect 3197 785 3203 1309
rect 3777 1309 3806 1334
rect 3174 760 3203 785
rect 3777 785 3783 1309
rect 3800 785 3806 1309
rect 3777 760 3806 785
rect 3174 754 3806 760
rect 3174 737 3228 754
rect 3752 737 3806 754
rect 3174 731 3806 737
rect 3872 1357 4504 1363
rect 3872 1340 3926 1357
rect 4450 1340 4504 1357
rect 3872 1334 4504 1340
rect 3872 1309 3901 1334
rect 3872 785 3878 1309
rect 3895 785 3901 1309
rect 4475 1309 4504 1334
rect 3872 760 3901 785
rect 4475 785 4481 1309
rect 4498 785 4504 1309
rect 4475 760 4504 785
rect 3872 754 4504 760
rect 3872 737 3926 754
rect 4450 737 4504 754
rect 3872 731 4504 737
rect 4570 1357 5202 1363
rect 4570 1340 4624 1357
rect 5148 1340 5202 1357
rect 4570 1334 5202 1340
rect 4570 1309 4599 1334
rect 4570 785 4576 1309
rect 4593 785 4599 1309
rect 5173 1309 5202 1334
rect 4570 760 4599 785
rect 5173 785 5179 1309
rect 5196 785 5202 1309
rect 5173 760 5202 785
rect 4570 754 5202 760
rect 4570 737 4624 754
rect 5148 737 5202 754
rect 4570 731 5202 737
rect -5202 659 -4570 665
rect -5202 642 -5148 659
rect -4624 642 -4570 659
rect -5202 636 -4570 642
rect -5202 611 -5173 636
rect -5202 87 -5196 611
rect -5179 87 -5173 611
rect -4599 611 -4570 636
rect -5202 62 -5173 87
rect -4599 87 -4593 611
rect -4576 87 -4570 611
rect -4599 62 -4570 87
rect -5202 56 -4570 62
rect -5202 39 -5148 56
rect -4624 39 -4570 56
rect -5202 33 -4570 39
rect -4504 659 -3872 665
rect -4504 642 -4450 659
rect -3926 642 -3872 659
rect -4504 636 -3872 642
rect -4504 611 -4475 636
rect -4504 87 -4498 611
rect -4481 87 -4475 611
rect -3901 611 -3872 636
rect -4504 62 -4475 87
rect -3901 87 -3895 611
rect -3878 87 -3872 611
rect -3901 62 -3872 87
rect -4504 56 -3872 62
rect -4504 39 -4450 56
rect -3926 39 -3872 56
rect -4504 33 -3872 39
rect -3806 659 -3174 665
rect -3806 642 -3752 659
rect -3228 642 -3174 659
rect -3806 636 -3174 642
rect -3806 611 -3777 636
rect -3806 87 -3800 611
rect -3783 87 -3777 611
rect -3203 611 -3174 636
rect -3806 62 -3777 87
rect -3203 87 -3197 611
rect -3180 87 -3174 611
rect -3203 62 -3174 87
rect -3806 56 -3174 62
rect -3806 39 -3752 56
rect -3228 39 -3174 56
rect -3806 33 -3174 39
rect -3108 659 -2476 665
rect -3108 642 -3054 659
rect -2530 642 -2476 659
rect -3108 636 -2476 642
rect -3108 611 -3079 636
rect -3108 87 -3102 611
rect -3085 87 -3079 611
rect -2505 611 -2476 636
rect -3108 62 -3079 87
rect -2505 87 -2499 611
rect -2482 87 -2476 611
rect -2505 62 -2476 87
rect -3108 56 -2476 62
rect -3108 39 -3054 56
rect -2530 39 -2476 56
rect -3108 33 -2476 39
rect -2410 659 -1778 665
rect -2410 642 -2356 659
rect -1832 642 -1778 659
rect -2410 636 -1778 642
rect -2410 611 -2381 636
rect -2410 87 -2404 611
rect -2387 87 -2381 611
rect -1807 611 -1778 636
rect -2410 62 -2381 87
rect -1807 87 -1801 611
rect -1784 87 -1778 611
rect -1807 62 -1778 87
rect -2410 56 -1778 62
rect -2410 39 -2356 56
rect -1832 39 -1778 56
rect -2410 33 -1778 39
rect -1712 659 -1080 665
rect -1712 642 -1658 659
rect -1134 642 -1080 659
rect -1712 636 -1080 642
rect -1712 611 -1683 636
rect -1712 87 -1706 611
rect -1689 87 -1683 611
rect -1109 611 -1080 636
rect -1712 62 -1683 87
rect -1109 87 -1103 611
rect -1086 87 -1080 611
rect -1109 62 -1080 87
rect -1712 56 -1080 62
rect -1712 39 -1658 56
rect -1134 39 -1080 56
rect -1712 33 -1080 39
rect -1014 659 -382 665
rect -1014 642 -960 659
rect -436 642 -382 659
rect -1014 636 -382 642
rect -1014 611 -985 636
rect -1014 87 -1008 611
rect -991 87 -985 611
rect -411 611 -382 636
rect -1014 62 -985 87
rect -411 87 -405 611
rect -388 87 -382 611
rect -411 62 -382 87
rect -1014 56 -382 62
rect -1014 39 -960 56
rect -436 39 -382 56
rect -1014 33 -382 39
rect -316 659 316 665
rect -316 642 -262 659
rect 262 642 316 659
rect -316 636 316 642
rect -316 611 -287 636
rect -316 87 -310 611
rect -293 87 -287 611
rect 287 611 316 636
rect -316 62 -287 87
rect 287 87 293 611
rect 310 87 316 611
rect 287 62 316 87
rect -316 56 316 62
rect -316 39 -262 56
rect 262 39 316 56
rect -316 33 316 39
rect 382 659 1014 665
rect 382 642 436 659
rect 960 642 1014 659
rect 382 636 1014 642
rect 382 611 411 636
rect 382 87 388 611
rect 405 87 411 611
rect 985 611 1014 636
rect 382 62 411 87
rect 985 87 991 611
rect 1008 87 1014 611
rect 985 62 1014 87
rect 382 56 1014 62
rect 382 39 436 56
rect 960 39 1014 56
rect 382 33 1014 39
rect 1080 659 1712 665
rect 1080 642 1134 659
rect 1658 642 1712 659
rect 1080 636 1712 642
rect 1080 611 1109 636
rect 1080 87 1086 611
rect 1103 87 1109 611
rect 1683 611 1712 636
rect 1080 62 1109 87
rect 1683 87 1689 611
rect 1706 87 1712 611
rect 1683 62 1712 87
rect 1080 56 1712 62
rect 1080 39 1134 56
rect 1658 39 1712 56
rect 1080 33 1712 39
rect 1778 659 2410 665
rect 1778 642 1832 659
rect 2356 642 2410 659
rect 1778 636 2410 642
rect 1778 611 1807 636
rect 1778 87 1784 611
rect 1801 87 1807 611
rect 2381 611 2410 636
rect 1778 62 1807 87
rect 2381 87 2387 611
rect 2404 87 2410 611
rect 2381 62 2410 87
rect 1778 56 2410 62
rect 1778 39 1832 56
rect 2356 39 2410 56
rect 1778 33 2410 39
rect 2476 659 3108 665
rect 2476 642 2530 659
rect 3054 642 3108 659
rect 2476 636 3108 642
rect 2476 611 2505 636
rect 2476 87 2482 611
rect 2499 87 2505 611
rect 3079 611 3108 636
rect 2476 62 2505 87
rect 3079 87 3085 611
rect 3102 87 3108 611
rect 3079 62 3108 87
rect 2476 56 3108 62
rect 2476 39 2530 56
rect 3054 39 3108 56
rect 2476 33 3108 39
rect 3174 659 3806 665
rect 3174 642 3228 659
rect 3752 642 3806 659
rect 3174 636 3806 642
rect 3174 611 3203 636
rect 3174 87 3180 611
rect 3197 87 3203 611
rect 3777 611 3806 636
rect 3174 62 3203 87
rect 3777 87 3783 611
rect 3800 87 3806 611
rect 3777 62 3806 87
rect 3174 56 3806 62
rect 3174 39 3228 56
rect 3752 39 3806 56
rect 3174 33 3806 39
rect 3872 659 4504 665
rect 3872 642 3926 659
rect 4450 642 4504 659
rect 3872 636 4504 642
rect 3872 611 3901 636
rect 3872 87 3878 611
rect 3895 87 3901 611
rect 4475 611 4504 636
rect 3872 62 3901 87
rect 4475 87 4481 611
rect 4498 87 4504 611
rect 4475 62 4504 87
rect 3872 56 4504 62
rect 3872 39 3926 56
rect 4450 39 4504 56
rect 3872 33 4504 39
rect 4570 659 5202 665
rect 4570 642 4624 659
rect 5148 642 5202 659
rect 4570 636 5202 642
rect 4570 611 4599 636
rect 4570 87 4576 611
rect 4593 87 4599 611
rect 5173 611 5202 636
rect 4570 62 4599 87
rect 5173 87 5179 611
rect 5196 87 5202 611
rect 5173 62 5202 87
rect 4570 56 5202 62
rect 4570 39 4624 56
rect 5148 39 5202 56
rect 4570 33 5202 39
rect -5202 -39 -4570 -33
rect -5202 -56 -5148 -39
rect -4624 -56 -4570 -39
rect -5202 -62 -4570 -56
rect -5202 -87 -5173 -62
rect -5202 -611 -5196 -87
rect -5179 -611 -5173 -87
rect -4599 -87 -4570 -62
rect -5202 -636 -5173 -611
rect -4599 -611 -4593 -87
rect -4576 -611 -4570 -87
rect -4599 -636 -4570 -611
rect -5202 -642 -4570 -636
rect -5202 -659 -5148 -642
rect -4624 -659 -4570 -642
rect -5202 -665 -4570 -659
rect -4504 -39 -3872 -33
rect -4504 -56 -4450 -39
rect -3926 -56 -3872 -39
rect -4504 -62 -3872 -56
rect -4504 -87 -4475 -62
rect -4504 -611 -4498 -87
rect -4481 -611 -4475 -87
rect -3901 -87 -3872 -62
rect -4504 -636 -4475 -611
rect -3901 -611 -3895 -87
rect -3878 -611 -3872 -87
rect -3901 -636 -3872 -611
rect -4504 -642 -3872 -636
rect -4504 -659 -4450 -642
rect -3926 -659 -3872 -642
rect -4504 -665 -3872 -659
rect -3806 -39 -3174 -33
rect -3806 -56 -3752 -39
rect -3228 -56 -3174 -39
rect -3806 -62 -3174 -56
rect -3806 -87 -3777 -62
rect -3806 -611 -3800 -87
rect -3783 -611 -3777 -87
rect -3203 -87 -3174 -62
rect -3806 -636 -3777 -611
rect -3203 -611 -3197 -87
rect -3180 -611 -3174 -87
rect -3203 -636 -3174 -611
rect -3806 -642 -3174 -636
rect -3806 -659 -3752 -642
rect -3228 -659 -3174 -642
rect -3806 -665 -3174 -659
rect -3108 -39 -2476 -33
rect -3108 -56 -3054 -39
rect -2530 -56 -2476 -39
rect -3108 -62 -2476 -56
rect -3108 -87 -3079 -62
rect -3108 -611 -3102 -87
rect -3085 -611 -3079 -87
rect -2505 -87 -2476 -62
rect -3108 -636 -3079 -611
rect -2505 -611 -2499 -87
rect -2482 -611 -2476 -87
rect -2505 -636 -2476 -611
rect -3108 -642 -2476 -636
rect -3108 -659 -3054 -642
rect -2530 -659 -2476 -642
rect -3108 -665 -2476 -659
rect -2410 -39 -1778 -33
rect -2410 -56 -2356 -39
rect -1832 -56 -1778 -39
rect -2410 -62 -1778 -56
rect -2410 -87 -2381 -62
rect -2410 -611 -2404 -87
rect -2387 -611 -2381 -87
rect -1807 -87 -1778 -62
rect -2410 -636 -2381 -611
rect -1807 -611 -1801 -87
rect -1784 -611 -1778 -87
rect -1807 -636 -1778 -611
rect -2410 -642 -1778 -636
rect -2410 -659 -2356 -642
rect -1832 -659 -1778 -642
rect -2410 -665 -1778 -659
rect -1712 -39 -1080 -33
rect -1712 -56 -1658 -39
rect -1134 -56 -1080 -39
rect -1712 -62 -1080 -56
rect -1712 -87 -1683 -62
rect -1712 -611 -1706 -87
rect -1689 -611 -1683 -87
rect -1109 -87 -1080 -62
rect -1712 -636 -1683 -611
rect -1109 -611 -1103 -87
rect -1086 -611 -1080 -87
rect -1109 -636 -1080 -611
rect -1712 -642 -1080 -636
rect -1712 -659 -1658 -642
rect -1134 -659 -1080 -642
rect -1712 -665 -1080 -659
rect -1014 -39 -382 -33
rect -1014 -56 -960 -39
rect -436 -56 -382 -39
rect -1014 -62 -382 -56
rect -1014 -87 -985 -62
rect -1014 -611 -1008 -87
rect -991 -611 -985 -87
rect -411 -87 -382 -62
rect -1014 -636 -985 -611
rect -411 -611 -405 -87
rect -388 -611 -382 -87
rect -411 -636 -382 -611
rect -1014 -642 -382 -636
rect -1014 -659 -960 -642
rect -436 -659 -382 -642
rect -1014 -665 -382 -659
rect -316 -39 316 -33
rect -316 -56 -262 -39
rect 262 -56 316 -39
rect -316 -62 316 -56
rect -316 -87 -287 -62
rect -316 -611 -310 -87
rect -293 -611 -287 -87
rect 287 -87 316 -62
rect -316 -636 -287 -611
rect 287 -611 293 -87
rect 310 -611 316 -87
rect 287 -636 316 -611
rect -316 -642 316 -636
rect -316 -659 -262 -642
rect 262 -659 316 -642
rect -316 -665 316 -659
rect 382 -39 1014 -33
rect 382 -56 436 -39
rect 960 -56 1014 -39
rect 382 -62 1014 -56
rect 382 -87 411 -62
rect 382 -611 388 -87
rect 405 -611 411 -87
rect 985 -87 1014 -62
rect 382 -636 411 -611
rect 985 -611 991 -87
rect 1008 -611 1014 -87
rect 985 -636 1014 -611
rect 382 -642 1014 -636
rect 382 -659 436 -642
rect 960 -659 1014 -642
rect 382 -665 1014 -659
rect 1080 -39 1712 -33
rect 1080 -56 1134 -39
rect 1658 -56 1712 -39
rect 1080 -62 1712 -56
rect 1080 -87 1109 -62
rect 1080 -611 1086 -87
rect 1103 -611 1109 -87
rect 1683 -87 1712 -62
rect 1080 -636 1109 -611
rect 1683 -611 1689 -87
rect 1706 -611 1712 -87
rect 1683 -636 1712 -611
rect 1080 -642 1712 -636
rect 1080 -659 1134 -642
rect 1658 -659 1712 -642
rect 1080 -665 1712 -659
rect 1778 -39 2410 -33
rect 1778 -56 1832 -39
rect 2356 -56 2410 -39
rect 1778 -62 2410 -56
rect 1778 -87 1807 -62
rect 1778 -611 1784 -87
rect 1801 -611 1807 -87
rect 2381 -87 2410 -62
rect 1778 -636 1807 -611
rect 2381 -611 2387 -87
rect 2404 -611 2410 -87
rect 2381 -636 2410 -611
rect 1778 -642 2410 -636
rect 1778 -659 1832 -642
rect 2356 -659 2410 -642
rect 1778 -665 2410 -659
rect 2476 -39 3108 -33
rect 2476 -56 2530 -39
rect 3054 -56 3108 -39
rect 2476 -62 3108 -56
rect 2476 -87 2505 -62
rect 2476 -611 2482 -87
rect 2499 -611 2505 -87
rect 3079 -87 3108 -62
rect 2476 -636 2505 -611
rect 3079 -611 3085 -87
rect 3102 -611 3108 -87
rect 3079 -636 3108 -611
rect 2476 -642 3108 -636
rect 2476 -659 2530 -642
rect 3054 -659 3108 -642
rect 2476 -665 3108 -659
rect 3174 -39 3806 -33
rect 3174 -56 3228 -39
rect 3752 -56 3806 -39
rect 3174 -62 3806 -56
rect 3174 -87 3203 -62
rect 3174 -611 3180 -87
rect 3197 -611 3203 -87
rect 3777 -87 3806 -62
rect 3174 -636 3203 -611
rect 3777 -611 3783 -87
rect 3800 -611 3806 -87
rect 3777 -636 3806 -611
rect 3174 -642 3806 -636
rect 3174 -659 3228 -642
rect 3752 -659 3806 -642
rect 3174 -665 3806 -659
rect 3872 -39 4504 -33
rect 3872 -56 3926 -39
rect 4450 -56 4504 -39
rect 3872 -62 4504 -56
rect 3872 -87 3901 -62
rect 3872 -611 3878 -87
rect 3895 -611 3901 -87
rect 4475 -87 4504 -62
rect 3872 -636 3901 -611
rect 4475 -611 4481 -87
rect 4498 -611 4504 -87
rect 4475 -636 4504 -611
rect 3872 -642 4504 -636
rect 3872 -659 3926 -642
rect 4450 -659 4504 -642
rect 3872 -665 4504 -659
rect 4570 -39 5202 -33
rect 4570 -56 4624 -39
rect 5148 -56 5202 -39
rect 4570 -62 5202 -56
rect 4570 -87 4599 -62
rect 4570 -611 4576 -87
rect 4593 -611 4599 -87
rect 5173 -87 5202 -62
rect 4570 -636 4599 -611
rect 5173 -611 5179 -87
rect 5196 -611 5202 -87
rect 5173 -636 5202 -611
rect 4570 -642 5202 -636
rect 4570 -659 4624 -642
rect 5148 -659 5202 -642
rect 4570 -665 5202 -659
rect -5202 -737 -4570 -731
rect -5202 -754 -5148 -737
rect -4624 -754 -4570 -737
rect -5202 -760 -4570 -754
rect -5202 -785 -5173 -760
rect -5202 -1309 -5196 -785
rect -5179 -1309 -5173 -785
rect -4599 -785 -4570 -760
rect -5202 -1334 -5173 -1309
rect -4599 -1309 -4593 -785
rect -4576 -1309 -4570 -785
rect -4599 -1334 -4570 -1309
rect -5202 -1340 -4570 -1334
rect -5202 -1357 -5148 -1340
rect -4624 -1357 -4570 -1340
rect -5202 -1363 -4570 -1357
rect -4504 -737 -3872 -731
rect -4504 -754 -4450 -737
rect -3926 -754 -3872 -737
rect -4504 -760 -3872 -754
rect -4504 -785 -4475 -760
rect -4504 -1309 -4498 -785
rect -4481 -1309 -4475 -785
rect -3901 -785 -3872 -760
rect -4504 -1334 -4475 -1309
rect -3901 -1309 -3895 -785
rect -3878 -1309 -3872 -785
rect -3901 -1334 -3872 -1309
rect -4504 -1340 -3872 -1334
rect -4504 -1357 -4450 -1340
rect -3926 -1357 -3872 -1340
rect -4504 -1363 -3872 -1357
rect -3806 -737 -3174 -731
rect -3806 -754 -3752 -737
rect -3228 -754 -3174 -737
rect -3806 -760 -3174 -754
rect -3806 -785 -3777 -760
rect -3806 -1309 -3800 -785
rect -3783 -1309 -3777 -785
rect -3203 -785 -3174 -760
rect -3806 -1334 -3777 -1309
rect -3203 -1309 -3197 -785
rect -3180 -1309 -3174 -785
rect -3203 -1334 -3174 -1309
rect -3806 -1340 -3174 -1334
rect -3806 -1357 -3752 -1340
rect -3228 -1357 -3174 -1340
rect -3806 -1363 -3174 -1357
rect -3108 -737 -2476 -731
rect -3108 -754 -3054 -737
rect -2530 -754 -2476 -737
rect -3108 -760 -2476 -754
rect -3108 -785 -3079 -760
rect -3108 -1309 -3102 -785
rect -3085 -1309 -3079 -785
rect -2505 -785 -2476 -760
rect -3108 -1334 -3079 -1309
rect -2505 -1309 -2499 -785
rect -2482 -1309 -2476 -785
rect -2505 -1334 -2476 -1309
rect -3108 -1340 -2476 -1334
rect -3108 -1357 -3054 -1340
rect -2530 -1357 -2476 -1340
rect -3108 -1363 -2476 -1357
rect -2410 -737 -1778 -731
rect -2410 -754 -2356 -737
rect -1832 -754 -1778 -737
rect -2410 -760 -1778 -754
rect -2410 -785 -2381 -760
rect -2410 -1309 -2404 -785
rect -2387 -1309 -2381 -785
rect -1807 -785 -1778 -760
rect -2410 -1334 -2381 -1309
rect -1807 -1309 -1801 -785
rect -1784 -1309 -1778 -785
rect -1807 -1334 -1778 -1309
rect -2410 -1340 -1778 -1334
rect -2410 -1357 -2356 -1340
rect -1832 -1357 -1778 -1340
rect -2410 -1363 -1778 -1357
rect -1712 -737 -1080 -731
rect -1712 -754 -1658 -737
rect -1134 -754 -1080 -737
rect -1712 -760 -1080 -754
rect -1712 -785 -1683 -760
rect -1712 -1309 -1706 -785
rect -1689 -1309 -1683 -785
rect -1109 -785 -1080 -760
rect -1712 -1334 -1683 -1309
rect -1109 -1309 -1103 -785
rect -1086 -1309 -1080 -785
rect -1109 -1334 -1080 -1309
rect -1712 -1340 -1080 -1334
rect -1712 -1357 -1658 -1340
rect -1134 -1357 -1080 -1340
rect -1712 -1363 -1080 -1357
rect -1014 -737 -382 -731
rect -1014 -754 -960 -737
rect -436 -754 -382 -737
rect -1014 -760 -382 -754
rect -1014 -785 -985 -760
rect -1014 -1309 -1008 -785
rect -991 -1309 -985 -785
rect -411 -785 -382 -760
rect -1014 -1334 -985 -1309
rect -411 -1309 -405 -785
rect -388 -1309 -382 -785
rect -411 -1334 -382 -1309
rect -1014 -1340 -382 -1334
rect -1014 -1357 -960 -1340
rect -436 -1357 -382 -1340
rect -1014 -1363 -382 -1357
rect -316 -737 316 -731
rect -316 -754 -262 -737
rect 262 -754 316 -737
rect -316 -760 316 -754
rect -316 -785 -287 -760
rect -316 -1309 -310 -785
rect -293 -1309 -287 -785
rect 287 -785 316 -760
rect -316 -1334 -287 -1309
rect 287 -1309 293 -785
rect 310 -1309 316 -785
rect 287 -1334 316 -1309
rect -316 -1340 316 -1334
rect -316 -1357 -262 -1340
rect 262 -1357 316 -1340
rect -316 -1363 316 -1357
rect 382 -737 1014 -731
rect 382 -754 436 -737
rect 960 -754 1014 -737
rect 382 -760 1014 -754
rect 382 -785 411 -760
rect 382 -1309 388 -785
rect 405 -1309 411 -785
rect 985 -785 1014 -760
rect 382 -1334 411 -1309
rect 985 -1309 991 -785
rect 1008 -1309 1014 -785
rect 985 -1334 1014 -1309
rect 382 -1340 1014 -1334
rect 382 -1357 436 -1340
rect 960 -1357 1014 -1340
rect 382 -1363 1014 -1357
rect 1080 -737 1712 -731
rect 1080 -754 1134 -737
rect 1658 -754 1712 -737
rect 1080 -760 1712 -754
rect 1080 -785 1109 -760
rect 1080 -1309 1086 -785
rect 1103 -1309 1109 -785
rect 1683 -785 1712 -760
rect 1080 -1334 1109 -1309
rect 1683 -1309 1689 -785
rect 1706 -1309 1712 -785
rect 1683 -1334 1712 -1309
rect 1080 -1340 1712 -1334
rect 1080 -1357 1134 -1340
rect 1658 -1357 1712 -1340
rect 1080 -1363 1712 -1357
rect 1778 -737 2410 -731
rect 1778 -754 1832 -737
rect 2356 -754 2410 -737
rect 1778 -760 2410 -754
rect 1778 -785 1807 -760
rect 1778 -1309 1784 -785
rect 1801 -1309 1807 -785
rect 2381 -785 2410 -760
rect 1778 -1334 1807 -1309
rect 2381 -1309 2387 -785
rect 2404 -1309 2410 -785
rect 2381 -1334 2410 -1309
rect 1778 -1340 2410 -1334
rect 1778 -1357 1832 -1340
rect 2356 -1357 2410 -1340
rect 1778 -1363 2410 -1357
rect 2476 -737 3108 -731
rect 2476 -754 2530 -737
rect 3054 -754 3108 -737
rect 2476 -760 3108 -754
rect 2476 -785 2505 -760
rect 2476 -1309 2482 -785
rect 2499 -1309 2505 -785
rect 3079 -785 3108 -760
rect 2476 -1334 2505 -1309
rect 3079 -1309 3085 -785
rect 3102 -1309 3108 -785
rect 3079 -1334 3108 -1309
rect 2476 -1340 3108 -1334
rect 2476 -1357 2530 -1340
rect 3054 -1357 3108 -1340
rect 2476 -1363 3108 -1357
rect 3174 -737 3806 -731
rect 3174 -754 3228 -737
rect 3752 -754 3806 -737
rect 3174 -760 3806 -754
rect 3174 -785 3203 -760
rect 3174 -1309 3180 -785
rect 3197 -1309 3203 -785
rect 3777 -785 3806 -760
rect 3174 -1334 3203 -1309
rect 3777 -1309 3783 -785
rect 3800 -1309 3806 -785
rect 3777 -1334 3806 -1309
rect 3174 -1340 3806 -1334
rect 3174 -1357 3228 -1340
rect 3752 -1357 3806 -1340
rect 3174 -1363 3806 -1357
rect 3872 -737 4504 -731
rect 3872 -754 3926 -737
rect 4450 -754 4504 -737
rect 3872 -760 4504 -754
rect 3872 -785 3901 -760
rect 3872 -1309 3878 -785
rect 3895 -1309 3901 -785
rect 4475 -785 4504 -760
rect 3872 -1334 3901 -1309
rect 4475 -1309 4481 -785
rect 4498 -1309 4504 -785
rect 4475 -1334 4504 -1309
rect 3872 -1340 4504 -1334
rect 3872 -1357 3926 -1340
rect 4450 -1357 4504 -1340
rect 3872 -1363 4504 -1357
rect 4570 -737 5202 -731
rect 4570 -754 4624 -737
rect 5148 -754 5202 -737
rect 4570 -760 5202 -754
rect 4570 -785 4599 -760
rect 4570 -1309 4576 -785
rect 4593 -1309 4599 -785
rect 5173 -785 5202 -760
rect 4570 -1334 4599 -1309
rect 5173 -1309 5179 -785
rect 5196 -1309 5202 -785
rect 5173 -1334 5202 -1309
rect 4570 -1340 5202 -1334
rect 4570 -1357 4624 -1340
rect 5148 -1357 5202 -1340
rect 4570 -1363 5202 -1357
<< mvpsubdiffcont >>
rect -5253 1445 5253 1462
rect -5301 -1414 -5284 1414
rect 5284 -1414 5301 1414
rect -5253 -1462 5253 -1445
<< mvnsubdiffcont >>
rect -5148 1340 -4624 1357
rect -5196 785 -5179 1309
rect -4593 785 -4576 1309
rect -5148 737 -4624 754
rect -4450 1340 -3926 1357
rect -4498 785 -4481 1309
rect -3895 785 -3878 1309
rect -4450 737 -3926 754
rect -3752 1340 -3228 1357
rect -3800 785 -3783 1309
rect -3197 785 -3180 1309
rect -3752 737 -3228 754
rect -3054 1340 -2530 1357
rect -3102 785 -3085 1309
rect -2499 785 -2482 1309
rect -3054 737 -2530 754
rect -2356 1340 -1832 1357
rect -2404 785 -2387 1309
rect -1801 785 -1784 1309
rect -2356 737 -1832 754
rect -1658 1340 -1134 1357
rect -1706 785 -1689 1309
rect -1103 785 -1086 1309
rect -1658 737 -1134 754
rect -960 1340 -436 1357
rect -1008 785 -991 1309
rect -405 785 -388 1309
rect -960 737 -436 754
rect -262 1340 262 1357
rect -310 785 -293 1309
rect 293 785 310 1309
rect -262 737 262 754
rect 436 1340 960 1357
rect 388 785 405 1309
rect 991 785 1008 1309
rect 436 737 960 754
rect 1134 1340 1658 1357
rect 1086 785 1103 1309
rect 1689 785 1706 1309
rect 1134 737 1658 754
rect 1832 1340 2356 1357
rect 1784 785 1801 1309
rect 2387 785 2404 1309
rect 1832 737 2356 754
rect 2530 1340 3054 1357
rect 2482 785 2499 1309
rect 3085 785 3102 1309
rect 2530 737 3054 754
rect 3228 1340 3752 1357
rect 3180 785 3197 1309
rect 3783 785 3800 1309
rect 3228 737 3752 754
rect 3926 1340 4450 1357
rect 3878 785 3895 1309
rect 4481 785 4498 1309
rect 3926 737 4450 754
rect 4624 1340 5148 1357
rect 4576 785 4593 1309
rect 5179 785 5196 1309
rect 4624 737 5148 754
rect -5148 642 -4624 659
rect -5196 87 -5179 611
rect -4593 87 -4576 611
rect -5148 39 -4624 56
rect -4450 642 -3926 659
rect -4498 87 -4481 611
rect -3895 87 -3878 611
rect -4450 39 -3926 56
rect -3752 642 -3228 659
rect -3800 87 -3783 611
rect -3197 87 -3180 611
rect -3752 39 -3228 56
rect -3054 642 -2530 659
rect -3102 87 -3085 611
rect -2499 87 -2482 611
rect -3054 39 -2530 56
rect -2356 642 -1832 659
rect -2404 87 -2387 611
rect -1801 87 -1784 611
rect -2356 39 -1832 56
rect -1658 642 -1134 659
rect -1706 87 -1689 611
rect -1103 87 -1086 611
rect -1658 39 -1134 56
rect -960 642 -436 659
rect -1008 87 -991 611
rect -405 87 -388 611
rect -960 39 -436 56
rect -262 642 262 659
rect -310 87 -293 611
rect 293 87 310 611
rect -262 39 262 56
rect 436 642 960 659
rect 388 87 405 611
rect 991 87 1008 611
rect 436 39 960 56
rect 1134 642 1658 659
rect 1086 87 1103 611
rect 1689 87 1706 611
rect 1134 39 1658 56
rect 1832 642 2356 659
rect 1784 87 1801 611
rect 2387 87 2404 611
rect 1832 39 2356 56
rect 2530 642 3054 659
rect 2482 87 2499 611
rect 3085 87 3102 611
rect 2530 39 3054 56
rect 3228 642 3752 659
rect 3180 87 3197 611
rect 3783 87 3800 611
rect 3228 39 3752 56
rect 3926 642 4450 659
rect 3878 87 3895 611
rect 4481 87 4498 611
rect 3926 39 4450 56
rect 4624 642 5148 659
rect 4576 87 4593 611
rect 5179 87 5196 611
rect 4624 39 5148 56
rect -5148 -56 -4624 -39
rect -5196 -611 -5179 -87
rect -4593 -611 -4576 -87
rect -5148 -659 -4624 -642
rect -4450 -56 -3926 -39
rect -4498 -611 -4481 -87
rect -3895 -611 -3878 -87
rect -4450 -659 -3926 -642
rect -3752 -56 -3228 -39
rect -3800 -611 -3783 -87
rect -3197 -611 -3180 -87
rect -3752 -659 -3228 -642
rect -3054 -56 -2530 -39
rect -3102 -611 -3085 -87
rect -2499 -611 -2482 -87
rect -3054 -659 -2530 -642
rect -2356 -56 -1832 -39
rect -2404 -611 -2387 -87
rect -1801 -611 -1784 -87
rect -2356 -659 -1832 -642
rect -1658 -56 -1134 -39
rect -1706 -611 -1689 -87
rect -1103 -611 -1086 -87
rect -1658 -659 -1134 -642
rect -960 -56 -436 -39
rect -1008 -611 -991 -87
rect -405 -611 -388 -87
rect -960 -659 -436 -642
rect -262 -56 262 -39
rect -310 -611 -293 -87
rect 293 -611 310 -87
rect -262 -659 262 -642
rect 436 -56 960 -39
rect 388 -611 405 -87
rect 991 -611 1008 -87
rect 436 -659 960 -642
rect 1134 -56 1658 -39
rect 1086 -611 1103 -87
rect 1689 -611 1706 -87
rect 1134 -659 1658 -642
rect 1832 -56 2356 -39
rect 1784 -611 1801 -87
rect 2387 -611 2404 -87
rect 1832 -659 2356 -642
rect 2530 -56 3054 -39
rect 2482 -611 2499 -87
rect 3085 -611 3102 -87
rect 2530 -659 3054 -642
rect 3228 -56 3752 -39
rect 3180 -611 3197 -87
rect 3783 -611 3800 -87
rect 3228 -659 3752 -642
rect 3926 -56 4450 -39
rect 3878 -611 3895 -87
rect 4481 -611 4498 -87
rect 3926 -659 4450 -642
rect 4624 -56 5148 -39
rect 4576 -611 4593 -87
rect 5179 -611 5196 -87
rect 4624 -659 5148 -642
rect -5148 -754 -4624 -737
rect -5196 -1309 -5179 -785
rect -4593 -1309 -4576 -785
rect -5148 -1357 -4624 -1340
rect -4450 -754 -3926 -737
rect -4498 -1309 -4481 -785
rect -3895 -1309 -3878 -785
rect -4450 -1357 -3926 -1340
rect -3752 -754 -3228 -737
rect -3800 -1309 -3783 -785
rect -3197 -1309 -3180 -785
rect -3752 -1357 -3228 -1340
rect -3054 -754 -2530 -737
rect -3102 -1309 -3085 -785
rect -2499 -1309 -2482 -785
rect -3054 -1357 -2530 -1340
rect -2356 -754 -1832 -737
rect -2404 -1309 -2387 -785
rect -1801 -1309 -1784 -785
rect -2356 -1357 -1832 -1340
rect -1658 -754 -1134 -737
rect -1706 -1309 -1689 -785
rect -1103 -1309 -1086 -785
rect -1658 -1357 -1134 -1340
rect -960 -754 -436 -737
rect -1008 -1309 -991 -785
rect -405 -1309 -388 -785
rect -960 -1357 -436 -1340
rect -262 -754 262 -737
rect -310 -1309 -293 -785
rect 293 -1309 310 -785
rect -262 -1357 262 -1340
rect 436 -754 960 -737
rect 388 -1309 405 -785
rect 991 -1309 1008 -785
rect 436 -1357 960 -1340
rect 1134 -754 1658 -737
rect 1086 -1309 1103 -785
rect 1689 -1309 1706 -785
rect 1134 -1357 1658 -1340
rect 1832 -754 2356 -737
rect 1784 -1309 1801 -785
rect 2387 -1309 2404 -785
rect 1832 -1357 2356 -1340
rect 2530 -754 3054 -737
rect 2482 -1309 2499 -785
rect 3085 -1309 3102 -785
rect 2530 -1357 3054 -1340
rect 3228 -754 3752 -737
rect 3180 -1309 3197 -785
rect 3783 -1309 3800 -785
rect 3228 -1357 3752 -1340
rect 3926 -754 4450 -737
rect 3878 -1309 3895 -785
rect 4481 -1309 4498 -785
rect 3926 -1357 4450 -1340
rect 4624 -754 5148 -737
rect 4576 -1309 4593 -785
rect 5179 -1309 5196 -785
rect 4624 -1357 5148 -1340
<< mvpdiode >>
rect -5136 1291 -4636 1297
rect -5136 803 -5130 1291
rect -4642 803 -4636 1291
rect -5136 797 -4636 803
rect -4438 1291 -3938 1297
rect -4438 803 -4432 1291
rect -3944 803 -3938 1291
rect -4438 797 -3938 803
rect -3740 1291 -3240 1297
rect -3740 803 -3734 1291
rect -3246 803 -3240 1291
rect -3740 797 -3240 803
rect -3042 1291 -2542 1297
rect -3042 803 -3036 1291
rect -2548 803 -2542 1291
rect -3042 797 -2542 803
rect -2344 1291 -1844 1297
rect -2344 803 -2338 1291
rect -1850 803 -1844 1291
rect -2344 797 -1844 803
rect -1646 1291 -1146 1297
rect -1646 803 -1640 1291
rect -1152 803 -1146 1291
rect -1646 797 -1146 803
rect -948 1291 -448 1297
rect -948 803 -942 1291
rect -454 803 -448 1291
rect -948 797 -448 803
rect -250 1291 250 1297
rect -250 803 -244 1291
rect 244 803 250 1291
rect -250 797 250 803
rect 448 1291 948 1297
rect 448 803 454 1291
rect 942 803 948 1291
rect 448 797 948 803
rect 1146 1291 1646 1297
rect 1146 803 1152 1291
rect 1640 803 1646 1291
rect 1146 797 1646 803
rect 1844 1291 2344 1297
rect 1844 803 1850 1291
rect 2338 803 2344 1291
rect 1844 797 2344 803
rect 2542 1291 3042 1297
rect 2542 803 2548 1291
rect 3036 803 3042 1291
rect 2542 797 3042 803
rect 3240 1291 3740 1297
rect 3240 803 3246 1291
rect 3734 803 3740 1291
rect 3240 797 3740 803
rect 3938 1291 4438 1297
rect 3938 803 3944 1291
rect 4432 803 4438 1291
rect 3938 797 4438 803
rect 4636 1291 5136 1297
rect 4636 803 4642 1291
rect 5130 803 5136 1291
rect 4636 797 5136 803
rect -5136 593 -4636 599
rect -5136 105 -5130 593
rect -4642 105 -4636 593
rect -5136 99 -4636 105
rect -4438 593 -3938 599
rect -4438 105 -4432 593
rect -3944 105 -3938 593
rect -4438 99 -3938 105
rect -3740 593 -3240 599
rect -3740 105 -3734 593
rect -3246 105 -3240 593
rect -3740 99 -3240 105
rect -3042 593 -2542 599
rect -3042 105 -3036 593
rect -2548 105 -2542 593
rect -3042 99 -2542 105
rect -2344 593 -1844 599
rect -2344 105 -2338 593
rect -1850 105 -1844 593
rect -2344 99 -1844 105
rect -1646 593 -1146 599
rect -1646 105 -1640 593
rect -1152 105 -1146 593
rect -1646 99 -1146 105
rect -948 593 -448 599
rect -948 105 -942 593
rect -454 105 -448 593
rect -948 99 -448 105
rect -250 593 250 599
rect -250 105 -244 593
rect 244 105 250 593
rect -250 99 250 105
rect 448 593 948 599
rect 448 105 454 593
rect 942 105 948 593
rect 448 99 948 105
rect 1146 593 1646 599
rect 1146 105 1152 593
rect 1640 105 1646 593
rect 1146 99 1646 105
rect 1844 593 2344 599
rect 1844 105 1850 593
rect 2338 105 2344 593
rect 1844 99 2344 105
rect 2542 593 3042 599
rect 2542 105 2548 593
rect 3036 105 3042 593
rect 2542 99 3042 105
rect 3240 593 3740 599
rect 3240 105 3246 593
rect 3734 105 3740 593
rect 3240 99 3740 105
rect 3938 593 4438 599
rect 3938 105 3944 593
rect 4432 105 4438 593
rect 3938 99 4438 105
rect 4636 593 5136 599
rect 4636 105 4642 593
rect 5130 105 5136 593
rect 4636 99 5136 105
rect -5136 -105 -4636 -99
rect -5136 -593 -5130 -105
rect -4642 -593 -4636 -105
rect -5136 -599 -4636 -593
rect -4438 -105 -3938 -99
rect -4438 -593 -4432 -105
rect -3944 -593 -3938 -105
rect -4438 -599 -3938 -593
rect -3740 -105 -3240 -99
rect -3740 -593 -3734 -105
rect -3246 -593 -3240 -105
rect -3740 -599 -3240 -593
rect -3042 -105 -2542 -99
rect -3042 -593 -3036 -105
rect -2548 -593 -2542 -105
rect -3042 -599 -2542 -593
rect -2344 -105 -1844 -99
rect -2344 -593 -2338 -105
rect -1850 -593 -1844 -105
rect -2344 -599 -1844 -593
rect -1646 -105 -1146 -99
rect -1646 -593 -1640 -105
rect -1152 -593 -1146 -105
rect -1646 -599 -1146 -593
rect -948 -105 -448 -99
rect -948 -593 -942 -105
rect -454 -593 -448 -105
rect -948 -599 -448 -593
rect -250 -105 250 -99
rect -250 -593 -244 -105
rect 244 -593 250 -105
rect -250 -599 250 -593
rect 448 -105 948 -99
rect 448 -593 454 -105
rect 942 -593 948 -105
rect 448 -599 948 -593
rect 1146 -105 1646 -99
rect 1146 -593 1152 -105
rect 1640 -593 1646 -105
rect 1146 -599 1646 -593
rect 1844 -105 2344 -99
rect 1844 -593 1850 -105
rect 2338 -593 2344 -105
rect 1844 -599 2344 -593
rect 2542 -105 3042 -99
rect 2542 -593 2548 -105
rect 3036 -593 3042 -105
rect 2542 -599 3042 -593
rect 3240 -105 3740 -99
rect 3240 -593 3246 -105
rect 3734 -593 3740 -105
rect 3240 -599 3740 -593
rect 3938 -105 4438 -99
rect 3938 -593 3944 -105
rect 4432 -593 4438 -105
rect 3938 -599 4438 -593
rect 4636 -105 5136 -99
rect 4636 -593 4642 -105
rect 5130 -593 5136 -105
rect 4636 -599 5136 -593
rect -5136 -803 -4636 -797
rect -5136 -1291 -5130 -803
rect -4642 -1291 -4636 -803
rect -5136 -1297 -4636 -1291
rect -4438 -803 -3938 -797
rect -4438 -1291 -4432 -803
rect -3944 -1291 -3938 -803
rect -4438 -1297 -3938 -1291
rect -3740 -803 -3240 -797
rect -3740 -1291 -3734 -803
rect -3246 -1291 -3240 -803
rect -3740 -1297 -3240 -1291
rect -3042 -803 -2542 -797
rect -3042 -1291 -3036 -803
rect -2548 -1291 -2542 -803
rect -3042 -1297 -2542 -1291
rect -2344 -803 -1844 -797
rect -2344 -1291 -2338 -803
rect -1850 -1291 -1844 -803
rect -2344 -1297 -1844 -1291
rect -1646 -803 -1146 -797
rect -1646 -1291 -1640 -803
rect -1152 -1291 -1146 -803
rect -1646 -1297 -1146 -1291
rect -948 -803 -448 -797
rect -948 -1291 -942 -803
rect -454 -1291 -448 -803
rect -948 -1297 -448 -1291
rect -250 -803 250 -797
rect -250 -1291 -244 -803
rect 244 -1291 250 -803
rect -250 -1297 250 -1291
rect 448 -803 948 -797
rect 448 -1291 454 -803
rect 942 -1291 948 -803
rect 448 -1297 948 -1291
rect 1146 -803 1646 -797
rect 1146 -1291 1152 -803
rect 1640 -1291 1646 -803
rect 1146 -1297 1646 -1291
rect 1844 -803 2344 -797
rect 1844 -1291 1850 -803
rect 2338 -1291 2344 -803
rect 1844 -1297 2344 -1291
rect 2542 -803 3042 -797
rect 2542 -1291 2548 -803
rect 3036 -1291 3042 -803
rect 2542 -1297 3042 -1291
rect 3240 -803 3740 -797
rect 3240 -1291 3246 -803
rect 3734 -1291 3740 -803
rect 3240 -1297 3740 -1291
rect 3938 -803 4438 -797
rect 3938 -1291 3944 -803
rect 4432 -1291 4438 -803
rect 3938 -1297 4438 -1291
rect 4636 -803 5136 -797
rect 4636 -1291 4642 -803
rect 5130 -1291 5136 -803
rect 4636 -1297 5136 -1291
<< mvpdiodec >>
rect -5130 803 -4642 1291
rect -4432 803 -3944 1291
rect -3734 803 -3246 1291
rect -3036 803 -2548 1291
rect -2338 803 -1850 1291
rect -1640 803 -1152 1291
rect -942 803 -454 1291
rect -244 803 244 1291
rect 454 803 942 1291
rect 1152 803 1640 1291
rect 1850 803 2338 1291
rect 2548 803 3036 1291
rect 3246 803 3734 1291
rect 3944 803 4432 1291
rect 4642 803 5130 1291
rect -5130 105 -4642 593
rect -4432 105 -3944 593
rect -3734 105 -3246 593
rect -3036 105 -2548 593
rect -2338 105 -1850 593
rect -1640 105 -1152 593
rect -942 105 -454 593
rect -244 105 244 593
rect 454 105 942 593
rect 1152 105 1640 593
rect 1850 105 2338 593
rect 2548 105 3036 593
rect 3246 105 3734 593
rect 3944 105 4432 593
rect 4642 105 5130 593
rect -5130 -593 -4642 -105
rect -4432 -593 -3944 -105
rect -3734 -593 -3246 -105
rect -3036 -593 -2548 -105
rect -2338 -593 -1850 -105
rect -1640 -593 -1152 -105
rect -942 -593 -454 -105
rect -244 -593 244 -105
rect 454 -593 942 -105
rect 1152 -593 1640 -105
rect 1850 -593 2338 -105
rect 2548 -593 3036 -105
rect 3246 -593 3734 -105
rect 3944 -593 4432 -105
rect 4642 -593 5130 -105
rect -5130 -1291 -4642 -803
rect -4432 -1291 -3944 -803
rect -3734 -1291 -3246 -803
rect -3036 -1291 -2548 -803
rect -2338 -1291 -1850 -803
rect -1640 -1291 -1152 -803
rect -942 -1291 -454 -803
rect -244 -1291 244 -803
rect 454 -1291 942 -803
rect 1152 -1291 1640 -803
rect 1850 -1291 2338 -803
rect 2548 -1291 3036 -803
rect 3246 -1291 3734 -803
rect 3944 -1291 4432 -803
rect 4642 -1291 5130 -803
<< locali >>
rect -5301 1445 -5253 1462
rect 5253 1445 5301 1462
rect -5301 1414 -5284 1445
rect 5284 1414 5301 1445
rect -5196 1340 -5148 1357
rect -4624 1340 -4576 1357
rect -5196 1309 -5179 1340
rect -4593 1309 -4576 1340
rect -5138 803 -5130 1291
rect -4642 803 -4634 1291
rect -5196 754 -5179 785
rect -4593 754 -4576 785
rect -5196 737 -5148 754
rect -4624 737 -4576 754
rect -4498 1340 -4450 1357
rect -3926 1340 -3878 1357
rect -4498 1309 -4481 1340
rect -3895 1309 -3878 1340
rect -4440 803 -4432 1291
rect -3944 803 -3936 1291
rect -4498 754 -4481 785
rect -3895 754 -3878 785
rect -4498 737 -4450 754
rect -3926 737 -3878 754
rect -3800 1340 -3752 1357
rect -3228 1340 -3180 1357
rect -3800 1309 -3783 1340
rect -3197 1309 -3180 1340
rect -3742 803 -3734 1291
rect -3246 803 -3238 1291
rect -3800 754 -3783 785
rect -3197 754 -3180 785
rect -3800 737 -3752 754
rect -3228 737 -3180 754
rect -3102 1340 -3054 1357
rect -2530 1340 -2482 1357
rect -3102 1309 -3085 1340
rect -2499 1309 -2482 1340
rect -3044 803 -3036 1291
rect -2548 803 -2540 1291
rect -3102 754 -3085 785
rect -2499 754 -2482 785
rect -3102 737 -3054 754
rect -2530 737 -2482 754
rect -2404 1340 -2356 1357
rect -1832 1340 -1784 1357
rect -2404 1309 -2387 1340
rect -1801 1309 -1784 1340
rect -2346 803 -2338 1291
rect -1850 803 -1842 1291
rect -2404 754 -2387 785
rect -1801 754 -1784 785
rect -2404 737 -2356 754
rect -1832 737 -1784 754
rect -1706 1340 -1658 1357
rect -1134 1340 -1086 1357
rect -1706 1309 -1689 1340
rect -1103 1309 -1086 1340
rect -1648 803 -1640 1291
rect -1152 803 -1144 1291
rect -1706 754 -1689 785
rect -1103 754 -1086 785
rect -1706 737 -1658 754
rect -1134 737 -1086 754
rect -1008 1340 -960 1357
rect -436 1340 -388 1357
rect -1008 1309 -991 1340
rect -405 1309 -388 1340
rect -950 803 -942 1291
rect -454 803 -446 1291
rect -1008 754 -991 785
rect -405 754 -388 785
rect -1008 737 -960 754
rect -436 737 -388 754
rect -310 1340 -262 1357
rect 262 1340 310 1357
rect -310 1309 -293 1340
rect 293 1309 310 1340
rect -252 803 -244 1291
rect 244 803 252 1291
rect -310 754 -293 785
rect 293 754 310 785
rect -310 737 -262 754
rect 262 737 310 754
rect 388 1340 436 1357
rect 960 1340 1008 1357
rect 388 1309 405 1340
rect 991 1309 1008 1340
rect 446 803 454 1291
rect 942 803 950 1291
rect 388 754 405 785
rect 991 754 1008 785
rect 388 737 436 754
rect 960 737 1008 754
rect 1086 1340 1134 1357
rect 1658 1340 1706 1357
rect 1086 1309 1103 1340
rect 1689 1309 1706 1340
rect 1144 803 1152 1291
rect 1640 803 1648 1291
rect 1086 754 1103 785
rect 1689 754 1706 785
rect 1086 737 1134 754
rect 1658 737 1706 754
rect 1784 1340 1832 1357
rect 2356 1340 2404 1357
rect 1784 1309 1801 1340
rect 2387 1309 2404 1340
rect 1842 803 1850 1291
rect 2338 803 2346 1291
rect 1784 754 1801 785
rect 2387 754 2404 785
rect 1784 737 1832 754
rect 2356 737 2404 754
rect 2482 1340 2530 1357
rect 3054 1340 3102 1357
rect 2482 1309 2499 1340
rect 3085 1309 3102 1340
rect 2540 803 2548 1291
rect 3036 803 3044 1291
rect 2482 754 2499 785
rect 3085 754 3102 785
rect 2482 737 2530 754
rect 3054 737 3102 754
rect 3180 1340 3228 1357
rect 3752 1340 3800 1357
rect 3180 1309 3197 1340
rect 3783 1309 3800 1340
rect 3238 803 3246 1291
rect 3734 803 3742 1291
rect 3180 754 3197 785
rect 3783 754 3800 785
rect 3180 737 3228 754
rect 3752 737 3800 754
rect 3878 1340 3926 1357
rect 4450 1340 4498 1357
rect 3878 1309 3895 1340
rect 4481 1309 4498 1340
rect 3936 803 3944 1291
rect 4432 803 4440 1291
rect 3878 754 3895 785
rect 4481 754 4498 785
rect 3878 737 3926 754
rect 4450 737 4498 754
rect 4576 1340 4624 1357
rect 5148 1340 5196 1357
rect 4576 1309 4593 1340
rect 5179 1309 5196 1340
rect 4634 803 4642 1291
rect 5130 803 5138 1291
rect 4576 754 4593 785
rect 5179 754 5196 785
rect 4576 737 4624 754
rect 5148 737 5196 754
rect -5196 642 -5148 659
rect -4624 642 -4576 659
rect -5196 611 -5179 642
rect -4593 611 -4576 642
rect -5138 105 -5130 593
rect -4642 105 -4634 593
rect -5196 56 -5179 87
rect -4593 56 -4576 87
rect -5196 39 -5148 56
rect -4624 39 -4576 56
rect -4498 642 -4450 659
rect -3926 642 -3878 659
rect -4498 611 -4481 642
rect -3895 611 -3878 642
rect -4440 105 -4432 593
rect -3944 105 -3936 593
rect -4498 56 -4481 87
rect -3895 56 -3878 87
rect -4498 39 -4450 56
rect -3926 39 -3878 56
rect -3800 642 -3752 659
rect -3228 642 -3180 659
rect -3800 611 -3783 642
rect -3197 611 -3180 642
rect -3742 105 -3734 593
rect -3246 105 -3238 593
rect -3800 56 -3783 87
rect -3197 56 -3180 87
rect -3800 39 -3752 56
rect -3228 39 -3180 56
rect -3102 642 -3054 659
rect -2530 642 -2482 659
rect -3102 611 -3085 642
rect -2499 611 -2482 642
rect -3044 105 -3036 593
rect -2548 105 -2540 593
rect -3102 56 -3085 87
rect -2499 56 -2482 87
rect -3102 39 -3054 56
rect -2530 39 -2482 56
rect -2404 642 -2356 659
rect -1832 642 -1784 659
rect -2404 611 -2387 642
rect -1801 611 -1784 642
rect -2346 105 -2338 593
rect -1850 105 -1842 593
rect -2404 56 -2387 87
rect -1801 56 -1784 87
rect -2404 39 -2356 56
rect -1832 39 -1784 56
rect -1706 642 -1658 659
rect -1134 642 -1086 659
rect -1706 611 -1689 642
rect -1103 611 -1086 642
rect -1648 105 -1640 593
rect -1152 105 -1144 593
rect -1706 56 -1689 87
rect -1103 56 -1086 87
rect -1706 39 -1658 56
rect -1134 39 -1086 56
rect -1008 642 -960 659
rect -436 642 -388 659
rect -1008 611 -991 642
rect -405 611 -388 642
rect -950 105 -942 593
rect -454 105 -446 593
rect -1008 56 -991 87
rect -405 56 -388 87
rect -1008 39 -960 56
rect -436 39 -388 56
rect -310 642 -262 659
rect 262 642 310 659
rect -310 611 -293 642
rect 293 611 310 642
rect -252 105 -244 593
rect 244 105 252 593
rect -310 56 -293 87
rect 293 56 310 87
rect -310 39 -262 56
rect 262 39 310 56
rect 388 642 436 659
rect 960 642 1008 659
rect 388 611 405 642
rect 991 611 1008 642
rect 446 105 454 593
rect 942 105 950 593
rect 388 56 405 87
rect 991 56 1008 87
rect 388 39 436 56
rect 960 39 1008 56
rect 1086 642 1134 659
rect 1658 642 1706 659
rect 1086 611 1103 642
rect 1689 611 1706 642
rect 1144 105 1152 593
rect 1640 105 1648 593
rect 1086 56 1103 87
rect 1689 56 1706 87
rect 1086 39 1134 56
rect 1658 39 1706 56
rect 1784 642 1832 659
rect 2356 642 2404 659
rect 1784 611 1801 642
rect 2387 611 2404 642
rect 1842 105 1850 593
rect 2338 105 2346 593
rect 1784 56 1801 87
rect 2387 56 2404 87
rect 1784 39 1832 56
rect 2356 39 2404 56
rect 2482 642 2530 659
rect 3054 642 3102 659
rect 2482 611 2499 642
rect 3085 611 3102 642
rect 2540 105 2548 593
rect 3036 105 3044 593
rect 2482 56 2499 87
rect 3085 56 3102 87
rect 2482 39 2530 56
rect 3054 39 3102 56
rect 3180 642 3228 659
rect 3752 642 3800 659
rect 3180 611 3197 642
rect 3783 611 3800 642
rect 3238 105 3246 593
rect 3734 105 3742 593
rect 3180 56 3197 87
rect 3783 56 3800 87
rect 3180 39 3228 56
rect 3752 39 3800 56
rect 3878 642 3926 659
rect 4450 642 4498 659
rect 3878 611 3895 642
rect 4481 611 4498 642
rect 3936 105 3944 593
rect 4432 105 4440 593
rect 3878 56 3895 87
rect 4481 56 4498 87
rect 3878 39 3926 56
rect 4450 39 4498 56
rect 4576 642 4624 659
rect 5148 642 5196 659
rect 4576 611 4593 642
rect 5179 611 5196 642
rect 4634 105 4642 593
rect 5130 105 5138 593
rect 4576 56 4593 87
rect 5179 56 5196 87
rect 4576 39 4624 56
rect 5148 39 5196 56
rect -5196 -56 -5148 -39
rect -4624 -56 -4576 -39
rect -5196 -87 -5179 -56
rect -4593 -87 -4576 -56
rect -5138 -593 -5130 -105
rect -4642 -593 -4634 -105
rect -5196 -642 -5179 -611
rect -4593 -642 -4576 -611
rect -5196 -659 -5148 -642
rect -4624 -659 -4576 -642
rect -4498 -56 -4450 -39
rect -3926 -56 -3878 -39
rect -4498 -87 -4481 -56
rect -3895 -87 -3878 -56
rect -4440 -593 -4432 -105
rect -3944 -593 -3936 -105
rect -4498 -642 -4481 -611
rect -3895 -642 -3878 -611
rect -4498 -659 -4450 -642
rect -3926 -659 -3878 -642
rect -3800 -56 -3752 -39
rect -3228 -56 -3180 -39
rect -3800 -87 -3783 -56
rect -3197 -87 -3180 -56
rect -3742 -593 -3734 -105
rect -3246 -593 -3238 -105
rect -3800 -642 -3783 -611
rect -3197 -642 -3180 -611
rect -3800 -659 -3752 -642
rect -3228 -659 -3180 -642
rect -3102 -56 -3054 -39
rect -2530 -56 -2482 -39
rect -3102 -87 -3085 -56
rect -2499 -87 -2482 -56
rect -3044 -593 -3036 -105
rect -2548 -593 -2540 -105
rect -3102 -642 -3085 -611
rect -2499 -642 -2482 -611
rect -3102 -659 -3054 -642
rect -2530 -659 -2482 -642
rect -2404 -56 -2356 -39
rect -1832 -56 -1784 -39
rect -2404 -87 -2387 -56
rect -1801 -87 -1784 -56
rect -2346 -593 -2338 -105
rect -1850 -593 -1842 -105
rect -2404 -642 -2387 -611
rect -1801 -642 -1784 -611
rect -2404 -659 -2356 -642
rect -1832 -659 -1784 -642
rect -1706 -56 -1658 -39
rect -1134 -56 -1086 -39
rect -1706 -87 -1689 -56
rect -1103 -87 -1086 -56
rect -1648 -593 -1640 -105
rect -1152 -593 -1144 -105
rect -1706 -642 -1689 -611
rect -1103 -642 -1086 -611
rect -1706 -659 -1658 -642
rect -1134 -659 -1086 -642
rect -1008 -56 -960 -39
rect -436 -56 -388 -39
rect -1008 -87 -991 -56
rect -405 -87 -388 -56
rect -950 -593 -942 -105
rect -454 -593 -446 -105
rect -1008 -642 -991 -611
rect -405 -642 -388 -611
rect -1008 -659 -960 -642
rect -436 -659 -388 -642
rect -310 -56 -262 -39
rect 262 -56 310 -39
rect -310 -87 -293 -56
rect 293 -87 310 -56
rect -252 -593 -244 -105
rect 244 -593 252 -105
rect -310 -642 -293 -611
rect 293 -642 310 -611
rect -310 -659 -262 -642
rect 262 -659 310 -642
rect 388 -56 436 -39
rect 960 -56 1008 -39
rect 388 -87 405 -56
rect 991 -87 1008 -56
rect 446 -593 454 -105
rect 942 -593 950 -105
rect 388 -642 405 -611
rect 991 -642 1008 -611
rect 388 -659 436 -642
rect 960 -659 1008 -642
rect 1086 -56 1134 -39
rect 1658 -56 1706 -39
rect 1086 -87 1103 -56
rect 1689 -87 1706 -56
rect 1144 -593 1152 -105
rect 1640 -593 1648 -105
rect 1086 -642 1103 -611
rect 1689 -642 1706 -611
rect 1086 -659 1134 -642
rect 1658 -659 1706 -642
rect 1784 -56 1832 -39
rect 2356 -56 2404 -39
rect 1784 -87 1801 -56
rect 2387 -87 2404 -56
rect 1842 -593 1850 -105
rect 2338 -593 2346 -105
rect 1784 -642 1801 -611
rect 2387 -642 2404 -611
rect 1784 -659 1832 -642
rect 2356 -659 2404 -642
rect 2482 -56 2530 -39
rect 3054 -56 3102 -39
rect 2482 -87 2499 -56
rect 3085 -87 3102 -56
rect 2540 -593 2548 -105
rect 3036 -593 3044 -105
rect 2482 -642 2499 -611
rect 3085 -642 3102 -611
rect 2482 -659 2530 -642
rect 3054 -659 3102 -642
rect 3180 -56 3228 -39
rect 3752 -56 3800 -39
rect 3180 -87 3197 -56
rect 3783 -87 3800 -56
rect 3238 -593 3246 -105
rect 3734 -593 3742 -105
rect 3180 -642 3197 -611
rect 3783 -642 3800 -611
rect 3180 -659 3228 -642
rect 3752 -659 3800 -642
rect 3878 -56 3926 -39
rect 4450 -56 4498 -39
rect 3878 -87 3895 -56
rect 4481 -87 4498 -56
rect 3936 -593 3944 -105
rect 4432 -593 4440 -105
rect 3878 -642 3895 -611
rect 4481 -642 4498 -611
rect 3878 -659 3926 -642
rect 4450 -659 4498 -642
rect 4576 -56 4624 -39
rect 5148 -56 5196 -39
rect 4576 -87 4593 -56
rect 5179 -87 5196 -56
rect 4634 -593 4642 -105
rect 5130 -593 5138 -105
rect 4576 -642 4593 -611
rect 5179 -642 5196 -611
rect 4576 -659 4624 -642
rect 5148 -659 5196 -642
rect -5196 -754 -5148 -737
rect -4624 -754 -4576 -737
rect -5196 -785 -5179 -754
rect -4593 -785 -4576 -754
rect -5138 -1291 -5130 -803
rect -4642 -1291 -4634 -803
rect -5196 -1340 -5179 -1309
rect -4593 -1340 -4576 -1309
rect -5196 -1357 -5148 -1340
rect -4624 -1357 -4576 -1340
rect -4498 -754 -4450 -737
rect -3926 -754 -3878 -737
rect -4498 -785 -4481 -754
rect -3895 -785 -3878 -754
rect -4440 -1291 -4432 -803
rect -3944 -1291 -3936 -803
rect -4498 -1340 -4481 -1309
rect -3895 -1340 -3878 -1309
rect -4498 -1357 -4450 -1340
rect -3926 -1357 -3878 -1340
rect -3800 -754 -3752 -737
rect -3228 -754 -3180 -737
rect -3800 -785 -3783 -754
rect -3197 -785 -3180 -754
rect -3742 -1291 -3734 -803
rect -3246 -1291 -3238 -803
rect -3800 -1340 -3783 -1309
rect -3197 -1340 -3180 -1309
rect -3800 -1357 -3752 -1340
rect -3228 -1357 -3180 -1340
rect -3102 -754 -3054 -737
rect -2530 -754 -2482 -737
rect -3102 -785 -3085 -754
rect -2499 -785 -2482 -754
rect -3044 -1291 -3036 -803
rect -2548 -1291 -2540 -803
rect -3102 -1340 -3085 -1309
rect -2499 -1340 -2482 -1309
rect -3102 -1357 -3054 -1340
rect -2530 -1357 -2482 -1340
rect -2404 -754 -2356 -737
rect -1832 -754 -1784 -737
rect -2404 -785 -2387 -754
rect -1801 -785 -1784 -754
rect -2346 -1291 -2338 -803
rect -1850 -1291 -1842 -803
rect -2404 -1340 -2387 -1309
rect -1801 -1340 -1784 -1309
rect -2404 -1357 -2356 -1340
rect -1832 -1357 -1784 -1340
rect -1706 -754 -1658 -737
rect -1134 -754 -1086 -737
rect -1706 -785 -1689 -754
rect -1103 -785 -1086 -754
rect -1648 -1291 -1640 -803
rect -1152 -1291 -1144 -803
rect -1706 -1340 -1689 -1309
rect -1103 -1340 -1086 -1309
rect -1706 -1357 -1658 -1340
rect -1134 -1357 -1086 -1340
rect -1008 -754 -960 -737
rect -436 -754 -388 -737
rect -1008 -785 -991 -754
rect -405 -785 -388 -754
rect -950 -1291 -942 -803
rect -454 -1291 -446 -803
rect -1008 -1340 -991 -1309
rect -405 -1340 -388 -1309
rect -1008 -1357 -960 -1340
rect -436 -1357 -388 -1340
rect -310 -754 -262 -737
rect 262 -754 310 -737
rect -310 -785 -293 -754
rect 293 -785 310 -754
rect -252 -1291 -244 -803
rect 244 -1291 252 -803
rect -310 -1340 -293 -1309
rect 293 -1340 310 -1309
rect -310 -1357 -262 -1340
rect 262 -1357 310 -1340
rect 388 -754 436 -737
rect 960 -754 1008 -737
rect 388 -785 405 -754
rect 991 -785 1008 -754
rect 446 -1291 454 -803
rect 942 -1291 950 -803
rect 388 -1340 405 -1309
rect 991 -1340 1008 -1309
rect 388 -1357 436 -1340
rect 960 -1357 1008 -1340
rect 1086 -754 1134 -737
rect 1658 -754 1706 -737
rect 1086 -785 1103 -754
rect 1689 -785 1706 -754
rect 1144 -1291 1152 -803
rect 1640 -1291 1648 -803
rect 1086 -1340 1103 -1309
rect 1689 -1340 1706 -1309
rect 1086 -1357 1134 -1340
rect 1658 -1357 1706 -1340
rect 1784 -754 1832 -737
rect 2356 -754 2404 -737
rect 1784 -785 1801 -754
rect 2387 -785 2404 -754
rect 1842 -1291 1850 -803
rect 2338 -1291 2346 -803
rect 1784 -1340 1801 -1309
rect 2387 -1340 2404 -1309
rect 1784 -1357 1832 -1340
rect 2356 -1357 2404 -1340
rect 2482 -754 2530 -737
rect 3054 -754 3102 -737
rect 2482 -785 2499 -754
rect 3085 -785 3102 -754
rect 2540 -1291 2548 -803
rect 3036 -1291 3044 -803
rect 2482 -1340 2499 -1309
rect 3085 -1340 3102 -1309
rect 2482 -1357 2530 -1340
rect 3054 -1357 3102 -1340
rect 3180 -754 3228 -737
rect 3752 -754 3800 -737
rect 3180 -785 3197 -754
rect 3783 -785 3800 -754
rect 3238 -1291 3246 -803
rect 3734 -1291 3742 -803
rect 3180 -1340 3197 -1309
rect 3783 -1340 3800 -1309
rect 3180 -1357 3228 -1340
rect 3752 -1357 3800 -1340
rect 3878 -754 3926 -737
rect 4450 -754 4498 -737
rect 3878 -785 3895 -754
rect 4481 -785 4498 -754
rect 3936 -1291 3944 -803
rect 4432 -1291 4440 -803
rect 3878 -1340 3895 -1309
rect 4481 -1340 4498 -1309
rect 3878 -1357 3926 -1340
rect 4450 -1357 4498 -1340
rect 4576 -754 4624 -737
rect 5148 -754 5196 -737
rect 4576 -785 4593 -754
rect 5179 -785 5196 -754
rect 4634 -1291 4642 -803
rect 5130 -1291 5138 -803
rect 4576 -1340 4593 -1309
rect 5179 -1340 5196 -1309
rect 4576 -1357 4624 -1340
rect 5148 -1357 5196 -1340
rect -5301 -1445 -5284 -1414
rect 5284 -1445 5301 -1414
rect -5301 -1462 -5253 -1445
rect 5253 -1462 5301 -1445
<< viali >>
rect -5130 803 -4642 1291
rect -4432 803 -3944 1291
rect -3734 803 -3246 1291
rect -3036 803 -2548 1291
rect -2338 803 -1850 1291
rect -1640 803 -1152 1291
rect -942 803 -454 1291
rect -244 803 244 1291
rect 454 803 942 1291
rect 1152 803 1640 1291
rect 1850 803 2338 1291
rect 2548 803 3036 1291
rect 3246 803 3734 1291
rect 3944 803 4432 1291
rect 4642 803 5130 1291
rect -5130 105 -4642 593
rect -4432 105 -3944 593
rect -3734 105 -3246 593
rect -3036 105 -2548 593
rect -2338 105 -1850 593
rect -1640 105 -1152 593
rect -942 105 -454 593
rect -244 105 244 593
rect 454 105 942 593
rect 1152 105 1640 593
rect 1850 105 2338 593
rect 2548 105 3036 593
rect 3246 105 3734 593
rect 3944 105 4432 593
rect 4642 105 5130 593
rect -5130 -593 -4642 -105
rect -4432 -593 -3944 -105
rect -3734 -593 -3246 -105
rect -3036 -593 -2548 -105
rect -2338 -593 -1850 -105
rect -1640 -593 -1152 -105
rect -942 -593 -454 -105
rect -244 -593 244 -105
rect 454 -593 942 -105
rect 1152 -593 1640 -105
rect 1850 -593 2338 -105
rect 2548 -593 3036 -105
rect 3246 -593 3734 -105
rect 3944 -593 4432 -105
rect 4642 -593 5130 -105
rect -5130 -1291 -4642 -803
rect -4432 -1291 -3944 -803
rect -3734 -1291 -3246 -803
rect -3036 -1291 -2548 -803
rect -2338 -1291 -1850 -803
rect -1640 -1291 -1152 -803
rect -942 -1291 -454 -803
rect -244 -1291 244 -803
rect 454 -1291 942 -803
rect 1152 -1291 1640 -803
rect 1850 -1291 2338 -803
rect 2548 -1291 3036 -803
rect 3246 -1291 3734 -803
rect 3944 -1291 4432 -803
rect 4642 -1291 5130 -803
<< metal1 >>
rect -5136 1291 -4636 1294
rect -5136 803 -5130 1291
rect -4642 803 -4636 1291
rect -5136 800 -4636 803
rect -4438 1291 -3938 1294
rect -4438 803 -4432 1291
rect -3944 803 -3938 1291
rect -4438 800 -3938 803
rect -3740 1291 -3240 1294
rect -3740 803 -3734 1291
rect -3246 803 -3240 1291
rect -3740 800 -3240 803
rect -3042 1291 -2542 1294
rect -3042 803 -3036 1291
rect -2548 803 -2542 1291
rect -3042 800 -2542 803
rect -2344 1291 -1844 1294
rect -2344 803 -2338 1291
rect -1850 803 -1844 1291
rect -2344 800 -1844 803
rect -1646 1291 -1146 1294
rect -1646 803 -1640 1291
rect -1152 803 -1146 1291
rect -1646 800 -1146 803
rect -948 1291 -448 1294
rect -948 803 -942 1291
rect -454 803 -448 1291
rect -948 800 -448 803
rect -250 1291 250 1294
rect -250 803 -244 1291
rect 244 803 250 1291
rect -250 800 250 803
rect 448 1291 948 1294
rect 448 803 454 1291
rect 942 803 948 1291
rect 448 800 948 803
rect 1146 1291 1646 1294
rect 1146 803 1152 1291
rect 1640 803 1646 1291
rect 1146 800 1646 803
rect 1844 1291 2344 1294
rect 1844 803 1850 1291
rect 2338 803 2344 1291
rect 1844 800 2344 803
rect 2542 1291 3042 1294
rect 2542 803 2548 1291
rect 3036 803 3042 1291
rect 2542 800 3042 803
rect 3240 1291 3740 1294
rect 3240 803 3246 1291
rect 3734 803 3740 1291
rect 3240 800 3740 803
rect 3938 1291 4438 1294
rect 3938 803 3944 1291
rect 4432 803 4438 1291
rect 3938 800 4438 803
rect 4636 1291 5136 1294
rect 4636 803 4642 1291
rect 5130 803 5136 1291
rect 4636 800 5136 803
rect -5136 593 -4636 596
rect -5136 105 -5130 593
rect -4642 105 -4636 593
rect -5136 102 -4636 105
rect -4438 593 -3938 596
rect -4438 105 -4432 593
rect -3944 105 -3938 593
rect -4438 102 -3938 105
rect -3740 593 -3240 596
rect -3740 105 -3734 593
rect -3246 105 -3240 593
rect -3740 102 -3240 105
rect -3042 593 -2542 596
rect -3042 105 -3036 593
rect -2548 105 -2542 593
rect -3042 102 -2542 105
rect -2344 593 -1844 596
rect -2344 105 -2338 593
rect -1850 105 -1844 593
rect -2344 102 -1844 105
rect -1646 593 -1146 596
rect -1646 105 -1640 593
rect -1152 105 -1146 593
rect -1646 102 -1146 105
rect -948 593 -448 596
rect -948 105 -942 593
rect -454 105 -448 593
rect -948 102 -448 105
rect -250 593 250 596
rect -250 105 -244 593
rect 244 105 250 593
rect -250 102 250 105
rect 448 593 948 596
rect 448 105 454 593
rect 942 105 948 593
rect 448 102 948 105
rect 1146 593 1646 596
rect 1146 105 1152 593
rect 1640 105 1646 593
rect 1146 102 1646 105
rect 1844 593 2344 596
rect 1844 105 1850 593
rect 2338 105 2344 593
rect 1844 102 2344 105
rect 2542 593 3042 596
rect 2542 105 2548 593
rect 3036 105 3042 593
rect 2542 102 3042 105
rect 3240 593 3740 596
rect 3240 105 3246 593
rect 3734 105 3740 593
rect 3240 102 3740 105
rect 3938 593 4438 596
rect 3938 105 3944 593
rect 4432 105 4438 593
rect 3938 102 4438 105
rect 4636 593 5136 596
rect 4636 105 4642 593
rect 5130 105 5136 593
rect 4636 102 5136 105
rect -5136 -105 -4636 -102
rect -5136 -593 -5130 -105
rect -4642 -593 -4636 -105
rect -5136 -596 -4636 -593
rect -4438 -105 -3938 -102
rect -4438 -593 -4432 -105
rect -3944 -593 -3938 -105
rect -4438 -596 -3938 -593
rect -3740 -105 -3240 -102
rect -3740 -593 -3734 -105
rect -3246 -593 -3240 -105
rect -3740 -596 -3240 -593
rect -3042 -105 -2542 -102
rect -3042 -593 -3036 -105
rect -2548 -593 -2542 -105
rect -3042 -596 -2542 -593
rect -2344 -105 -1844 -102
rect -2344 -593 -2338 -105
rect -1850 -593 -1844 -105
rect -2344 -596 -1844 -593
rect -1646 -105 -1146 -102
rect -1646 -593 -1640 -105
rect -1152 -593 -1146 -105
rect -1646 -596 -1146 -593
rect -948 -105 -448 -102
rect -948 -593 -942 -105
rect -454 -593 -448 -105
rect -948 -596 -448 -593
rect -250 -105 250 -102
rect -250 -593 -244 -105
rect 244 -593 250 -105
rect -250 -596 250 -593
rect 448 -105 948 -102
rect 448 -593 454 -105
rect 942 -593 948 -105
rect 448 -596 948 -593
rect 1146 -105 1646 -102
rect 1146 -593 1152 -105
rect 1640 -593 1646 -105
rect 1146 -596 1646 -593
rect 1844 -105 2344 -102
rect 1844 -593 1850 -105
rect 2338 -593 2344 -105
rect 1844 -596 2344 -593
rect 2542 -105 3042 -102
rect 2542 -593 2548 -105
rect 3036 -593 3042 -105
rect 2542 -596 3042 -593
rect 3240 -105 3740 -102
rect 3240 -593 3246 -105
rect 3734 -593 3740 -105
rect 3240 -596 3740 -593
rect 3938 -105 4438 -102
rect 3938 -593 3944 -105
rect 4432 -593 4438 -105
rect 3938 -596 4438 -593
rect 4636 -105 5136 -102
rect 4636 -593 4642 -105
rect 5130 -593 5136 -105
rect 4636 -596 5136 -593
rect -5136 -803 -4636 -800
rect -5136 -1291 -5130 -803
rect -4642 -1291 -4636 -803
rect -5136 -1294 -4636 -1291
rect -4438 -803 -3938 -800
rect -4438 -1291 -4432 -803
rect -3944 -1291 -3938 -803
rect -4438 -1294 -3938 -1291
rect -3740 -803 -3240 -800
rect -3740 -1291 -3734 -803
rect -3246 -1291 -3240 -803
rect -3740 -1294 -3240 -1291
rect -3042 -803 -2542 -800
rect -3042 -1291 -3036 -803
rect -2548 -1291 -2542 -803
rect -3042 -1294 -2542 -1291
rect -2344 -803 -1844 -800
rect -2344 -1291 -2338 -803
rect -1850 -1291 -1844 -803
rect -2344 -1294 -1844 -1291
rect -1646 -803 -1146 -800
rect -1646 -1291 -1640 -803
rect -1152 -1291 -1146 -803
rect -1646 -1294 -1146 -1291
rect -948 -803 -448 -800
rect -948 -1291 -942 -803
rect -454 -1291 -448 -803
rect -948 -1294 -448 -1291
rect -250 -803 250 -800
rect -250 -1291 -244 -803
rect 244 -1291 250 -803
rect -250 -1294 250 -1291
rect 448 -803 948 -800
rect 448 -1291 454 -803
rect 942 -1291 948 -803
rect 448 -1294 948 -1291
rect 1146 -803 1646 -800
rect 1146 -1291 1152 -803
rect 1640 -1291 1646 -803
rect 1146 -1294 1646 -1291
rect 1844 -803 2344 -800
rect 1844 -1291 1850 -803
rect 2338 -1291 2344 -803
rect 1844 -1294 2344 -1291
rect 2542 -803 3042 -800
rect 2542 -1291 2548 -803
rect 3036 -1291 3042 -803
rect 2542 -1294 3042 -1291
rect 3240 -803 3740 -800
rect 3240 -1291 3246 -803
rect 3734 -1291 3740 -803
rect 3240 -1294 3740 -1291
rect 3938 -803 4438 -800
rect 3938 -1291 3944 -803
rect 4432 -1291 4438 -803
rect 3938 -1294 4438 -1291
rect 4636 -803 5136 -800
rect 4636 -1291 4642 -803
rect 5130 -1291 5136 -803
rect 4636 -1294 5136 -1291
<< properties >>
string FIXED_BBOX 4584 745 5187 1348
string gencell sky130_fd_pr__diode_pd2nw_11v0
string library sky130
string parameters w 5 l 5 area 25.0 peri 20.0 nx 15 ny 4 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 0 compatible {sky130_fd_pr__diode_pd2nw_05v5 sky130_fd_pr__diode_pd2nw_05v5_lvt  sky130_fd_pr__diode_pd2nw_05v5_hvt sky130_fd_pr__diode_pd2nw_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
