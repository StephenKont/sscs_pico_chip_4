magic
tech sky130A
timestamp 1665674841
<< nwell >>
rect -698 -2792 698 2792
<< pwell >>
rect -788 2792 788 2882
rect -788 -2792 -698 2792
rect 698 -2792 788 2792
rect -788 -2882 788 -2792
<< mvpsubdiff >>
rect -770 2858 770 2864
rect -770 2841 -716 2858
rect 716 2841 770 2858
rect -770 2835 770 2841
rect -770 2810 -741 2835
rect -770 -2810 -764 2810
rect -747 -2810 -741 2810
rect 741 2810 770 2835
rect -770 -2835 -741 -2810
rect 741 -2810 747 2810
rect 764 -2810 770 2810
rect 741 -2835 770 -2810
rect -770 -2841 770 -2835
rect -770 -2858 -716 -2841
rect 716 -2858 770 -2841
rect -770 -2864 770 -2858
<< mvnsubdiff >>
rect -665 2753 -33 2759
rect -665 2736 -611 2753
rect -87 2736 -33 2753
rect -665 2730 -33 2736
rect -665 2705 -636 2730
rect -665 2181 -659 2705
rect -642 2181 -636 2705
rect -62 2705 -33 2730
rect -665 2156 -636 2181
rect -62 2181 -56 2705
rect -39 2181 -33 2705
rect -62 2156 -33 2181
rect -665 2150 -33 2156
rect -665 2133 -611 2150
rect -87 2133 -33 2150
rect -665 2127 -33 2133
rect 33 2753 665 2759
rect 33 2736 87 2753
rect 611 2736 665 2753
rect 33 2730 665 2736
rect 33 2705 62 2730
rect 33 2181 39 2705
rect 56 2181 62 2705
rect 636 2705 665 2730
rect 33 2156 62 2181
rect 636 2181 642 2705
rect 659 2181 665 2705
rect 636 2156 665 2181
rect 33 2150 665 2156
rect 33 2133 87 2150
rect 611 2133 665 2150
rect 33 2127 665 2133
rect -665 2055 -33 2061
rect -665 2038 -611 2055
rect -87 2038 -33 2055
rect -665 2032 -33 2038
rect -665 2007 -636 2032
rect -665 1483 -659 2007
rect -642 1483 -636 2007
rect -62 2007 -33 2032
rect -665 1458 -636 1483
rect -62 1483 -56 2007
rect -39 1483 -33 2007
rect -62 1458 -33 1483
rect -665 1452 -33 1458
rect -665 1435 -611 1452
rect -87 1435 -33 1452
rect -665 1429 -33 1435
rect 33 2055 665 2061
rect 33 2038 87 2055
rect 611 2038 665 2055
rect 33 2032 665 2038
rect 33 2007 62 2032
rect 33 1483 39 2007
rect 56 1483 62 2007
rect 636 2007 665 2032
rect 33 1458 62 1483
rect 636 1483 642 2007
rect 659 1483 665 2007
rect 636 1458 665 1483
rect 33 1452 665 1458
rect 33 1435 87 1452
rect 611 1435 665 1452
rect 33 1429 665 1435
rect -665 1357 -33 1363
rect -665 1340 -611 1357
rect -87 1340 -33 1357
rect -665 1334 -33 1340
rect -665 1309 -636 1334
rect -665 785 -659 1309
rect -642 785 -636 1309
rect -62 1309 -33 1334
rect -665 760 -636 785
rect -62 785 -56 1309
rect -39 785 -33 1309
rect -62 760 -33 785
rect -665 754 -33 760
rect -665 737 -611 754
rect -87 737 -33 754
rect -665 731 -33 737
rect 33 1357 665 1363
rect 33 1340 87 1357
rect 611 1340 665 1357
rect 33 1334 665 1340
rect 33 1309 62 1334
rect 33 785 39 1309
rect 56 785 62 1309
rect 636 1309 665 1334
rect 33 760 62 785
rect 636 785 642 1309
rect 659 785 665 1309
rect 636 760 665 785
rect 33 754 665 760
rect 33 737 87 754
rect 611 737 665 754
rect 33 731 665 737
rect -665 659 -33 665
rect -665 642 -611 659
rect -87 642 -33 659
rect -665 636 -33 642
rect -665 611 -636 636
rect -665 87 -659 611
rect -642 87 -636 611
rect -62 611 -33 636
rect -665 62 -636 87
rect -62 87 -56 611
rect -39 87 -33 611
rect -62 62 -33 87
rect -665 56 -33 62
rect -665 39 -611 56
rect -87 39 -33 56
rect -665 33 -33 39
rect 33 659 665 665
rect 33 642 87 659
rect 611 642 665 659
rect 33 636 665 642
rect 33 611 62 636
rect 33 87 39 611
rect 56 87 62 611
rect 636 611 665 636
rect 33 62 62 87
rect 636 87 642 611
rect 659 87 665 611
rect 636 62 665 87
rect 33 56 665 62
rect 33 39 87 56
rect 611 39 665 56
rect 33 33 665 39
rect -665 -39 -33 -33
rect -665 -56 -611 -39
rect -87 -56 -33 -39
rect -665 -62 -33 -56
rect -665 -87 -636 -62
rect -665 -611 -659 -87
rect -642 -611 -636 -87
rect -62 -87 -33 -62
rect -665 -636 -636 -611
rect -62 -611 -56 -87
rect -39 -611 -33 -87
rect -62 -636 -33 -611
rect -665 -642 -33 -636
rect -665 -659 -611 -642
rect -87 -659 -33 -642
rect -665 -665 -33 -659
rect 33 -39 665 -33
rect 33 -56 87 -39
rect 611 -56 665 -39
rect 33 -62 665 -56
rect 33 -87 62 -62
rect 33 -611 39 -87
rect 56 -611 62 -87
rect 636 -87 665 -62
rect 33 -636 62 -611
rect 636 -611 642 -87
rect 659 -611 665 -87
rect 636 -636 665 -611
rect 33 -642 665 -636
rect 33 -659 87 -642
rect 611 -659 665 -642
rect 33 -665 665 -659
rect -665 -737 -33 -731
rect -665 -754 -611 -737
rect -87 -754 -33 -737
rect -665 -760 -33 -754
rect -665 -785 -636 -760
rect -665 -1309 -659 -785
rect -642 -1309 -636 -785
rect -62 -785 -33 -760
rect -665 -1334 -636 -1309
rect -62 -1309 -56 -785
rect -39 -1309 -33 -785
rect -62 -1334 -33 -1309
rect -665 -1340 -33 -1334
rect -665 -1357 -611 -1340
rect -87 -1357 -33 -1340
rect -665 -1363 -33 -1357
rect 33 -737 665 -731
rect 33 -754 87 -737
rect 611 -754 665 -737
rect 33 -760 665 -754
rect 33 -785 62 -760
rect 33 -1309 39 -785
rect 56 -1309 62 -785
rect 636 -785 665 -760
rect 33 -1334 62 -1309
rect 636 -1309 642 -785
rect 659 -1309 665 -785
rect 636 -1334 665 -1309
rect 33 -1340 665 -1334
rect 33 -1357 87 -1340
rect 611 -1357 665 -1340
rect 33 -1363 665 -1357
rect -665 -1435 -33 -1429
rect -665 -1452 -611 -1435
rect -87 -1452 -33 -1435
rect -665 -1458 -33 -1452
rect -665 -1483 -636 -1458
rect -665 -2007 -659 -1483
rect -642 -2007 -636 -1483
rect -62 -1483 -33 -1458
rect -665 -2032 -636 -2007
rect -62 -2007 -56 -1483
rect -39 -2007 -33 -1483
rect -62 -2032 -33 -2007
rect -665 -2038 -33 -2032
rect -665 -2055 -611 -2038
rect -87 -2055 -33 -2038
rect -665 -2061 -33 -2055
rect 33 -1435 665 -1429
rect 33 -1452 87 -1435
rect 611 -1452 665 -1435
rect 33 -1458 665 -1452
rect 33 -1483 62 -1458
rect 33 -2007 39 -1483
rect 56 -2007 62 -1483
rect 636 -1483 665 -1458
rect 33 -2032 62 -2007
rect 636 -2007 642 -1483
rect 659 -2007 665 -1483
rect 636 -2032 665 -2007
rect 33 -2038 665 -2032
rect 33 -2055 87 -2038
rect 611 -2055 665 -2038
rect 33 -2061 665 -2055
rect -665 -2133 -33 -2127
rect -665 -2150 -611 -2133
rect -87 -2150 -33 -2133
rect -665 -2156 -33 -2150
rect -665 -2181 -636 -2156
rect -665 -2705 -659 -2181
rect -642 -2705 -636 -2181
rect -62 -2181 -33 -2156
rect -665 -2730 -636 -2705
rect -62 -2705 -56 -2181
rect -39 -2705 -33 -2181
rect -62 -2730 -33 -2705
rect -665 -2736 -33 -2730
rect -665 -2753 -611 -2736
rect -87 -2753 -33 -2736
rect -665 -2759 -33 -2753
rect 33 -2133 665 -2127
rect 33 -2150 87 -2133
rect 611 -2150 665 -2133
rect 33 -2156 665 -2150
rect 33 -2181 62 -2156
rect 33 -2705 39 -2181
rect 56 -2705 62 -2181
rect 636 -2181 665 -2156
rect 33 -2730 62 -2705
rect 636 -2705 642 -2181
rect 659 -2705 665 -2181
rect 636 -2730 665 -2705
rect 33 -2736 665 -2730
rect 33 -2753 87 -2736
rect 611 -2753 665 -2736
rect 33 -2759 665 -2753
<< mvpsubdiffcont >>
rect -716 2841 716 2858
rect -764 -2810 -747 2810
rect 747 -2810 764 2810
rect -716 -2858 716 -2841
<< mvnsubdiffcont >>
rect -611 2736 -87 2753
rect -659 2181 -642 2705
rect -56 2181 -39 2705
rect -611 2133 -87 2150
rect 87 2736 611 2753
rect 39 2181 56 2705
rect 642 2181 659 2705
rect 87 2133 611 2150
rect -611 2038 -87 2055
rect -659 1483 -642 2007
rect -56 1483 -39 2007
rect -611 1435 -87 1452
rect 87 2038 611 2055
rect 39 1483 56 2007
rect 642 1483 659 2007
rect 87 1435 611 1452
rect -611 1340 -87 1357
rect -659 785 -642 1309
rect -56 785 -39 1309
rect -611 737 -87 754
rect 87 1340 611 1357
rect 39 785 56 1309
rect 642 785 659 1309
rect 87 737 611 754
rect -611 642 -87 659
rect -659 87 -642 611
rect -56 87 -39 611
rect -611 39 -87 56
rect 87 642 611 659
rect 39 87 56 611
rect 642 87 659 611
rect 87 39 611 56
rect -611 -56 -87 -39
rect -659 -611 -642 -87
rect -56 -611 -39 -87
rect -611 -659 -87 -642
rect 87 -56 611 -39
rect 39 -611 56 -87
rect 642 -611 659 -87
rect 87 -659 611 -642
rect -611 -754 -87 -737
rect -659 -1309 -642 -785
rect -56 -1309 -39 -785
rect -611 -1357 -87 -1340
rect 87 -754 611 -737
rect 39 -1309 56 -785
rect 642 -1309 659 -785
rect 87 -1357 611 -1340
rect -611 -1452 -87 -1435
rect -659 -2007 -642 -1483
rect -56 -2007 -39 -1483
rect -611 -2055 -87 -2038
rect 87 -1452 611 -1435
rect 39 -2007 56 -1483
rect 642 -2007 659 -1483
rect 87 -2055 611 -2038
rect -611 -2150 -87 -2133
rect -659 -2705 -642 -2181
rect -56 -2705 -39 -2181
rect -611 -2753 -87 -2736
rect 87 -2150 611 -2133
rect 39 -2705 56 -2181
rect 642 -2705 659 -2181
rect 87 -2753 611 -2736
<< mvpdiode >>
rect -599 2687 -99 2693
rect -599 2199 -593 2687
rect -105 2199 -99 2687
rect -599 2193 -99 2199
rect 99 2687 599 2693
rect 99 2199 105 2687
rect 593 2199 599 2687
rect 99 2193 599 2199
rect -599 1989 -99 1995
rect -599 1501 -593 1989
rect -105 1501 -99 1989
rect -599 1495 -99 1501
rect 99 1989 599 1995
rect 99 1501 105 1989
rect 593 1501 599 1989
rect 99 1495 599 1501
rect -599 1291 -99 1297
rect -599 803 -593 1291
rect -105 803 -99 1291
rect -599 797 -99 803
rect 99 1291 599 1297
rect 99 803 105 1291
rect 593 803 599 1291
rect 99 797 599 803
rect -599 593 -99 599
rect -599 105 -593 593
rect -105 105 -99 593
rect -599 99 -99 105
rect 99 593 599 599
rect 99 105 105 593
rect 593 105 599 593
rect 99 99 599 105
rect -599 -105 -99 -99
rect -599 -593 -593 -105
rect -105 -593 -99 -105
rect -599 -599 -99 -593
rect 99 -105 599 -99
rect 99 -593 105 -105
rect 593 -593 599 -105
rect 99 -599 599 -593
rect -599 -803 -99 -797
rect -599 -1291 -593 -803
rect -105 -1291 -99 -803
rect -599 -1297 -99 -1291
rect 99 -803 599 -797
rect 99 -1291 105 -803
rect 593 -1291 599 -803
rect 99 -1297 599 -1291
rect -599 -1501 -99 -1495
rect -599 -1989 -593 -1501
rect -105 -1989 -99 -1501
rect -599 -1995 -99 -1989
rect 99 -1501 599 -1495
rect 99 -1989 105 -1501
rect 593 -1989 599 -1501
rect 99 -1995 599 -1989
rect -599 -2199 -99 -2193
rect -599 -2687 -593 -2199
rect -105 -2687 -99 -2199
rect -599 -2693 -99 -2687
rect 99 -2199 599 -2193
rect 99 -2687 105 -2199
rect 593 -2687 599 -2199
rect 99 -2693 599 -2687
<< mvpdiodec >>
rect -593 2199 -105 2687
rect 105 2199 593 2687
rect -593 1501 -105 1989
rect 105 1501 593 1989
rect -593 803 -105 1291
rect 105 803 593 1291
rect -593 105 -105 593
rect 105 105 593 593
rect -593 -593 -105 -105
rect 105 -593 593 -105
rect -593 -1291 -105 -803
rect 105 -1291 593 -803
rect -593 -1989 -105 -1501
rect 105 -1989 593 -1501
rect -593 -2687 -105 -2199
rect 105 -2687 593 -2199
<< locali >>
rect -764 2841 -716 2858
rect 716 2841 764 2858
rect -764 2810 -747 2841
rect 747 2810 764 2841
rect -659 2736 -611 2753
rect -87 2736 -39 2753
rect -659 2705 -642 2736
rect -56 2705 -39 2736
rect -601 2199 -593 2687
rect -105 2199 -97 2687
rect -659 2150 -642 2181
rect -56 2150 -39 2181
rect -659 2133 -611 2150
rect -87 2133 -39 2150
rect 39 2736 87 2753
rect 611 2736 659 2753
rect 39 2705 56 2736
rect 642 2705 659 2736
rect 97 2199 105 2687
rect 593 2199 601 2687
rect 39 2150 56 2181
rect 642 2150 659 2181
rect 39 2133 87 2150
rect 611 2133 659 2150
rect -659 2038 -611 2055
rect -87 2038 -39 2055
rect -659 2007 -642 2038
rect -56 2007 -39 2038
rect -601 1501 -593 1989
rect -105 1501 -97 1989
rect -659 1452 -642 1483
rect -56 1452 -39 1483
rect -659 1435 -611 1452
rect -87 1435 -39 1452
rect 39 2038 87 2055
rect 611 2038 659 2055
rect 39 2007 56 2038
rect 642 2007 659 2038
rect 97 1501 105 1989
rect 593 1501 601 1989
rect 39 1452 56 1483
rect 642 1452 659 1483
rect 39 1435 87 1452
rect 611 1435 659 1452
rect -659 1340 -611 1357
rect -87 1340 -39 1357
rect -659 1309 -642 1340
rect -56 1309 -39 1340
rect -601 803 -593 1291
rect -105 803 -97 1291
rect -659 754 -642 785
rect -56 754 -39 785
rect -659 737 -611 754
rect -87 737 -39 754
rect 39 1340 87 1357
rect 611 1340 659 1357
rect 39 1309 56 1340
rect 642 1309 659 1340
rect 97 803 105 1291
rect 593 803 601 1291
rect 39 754 56 785
rect 642 754 659 785
rect 39 737 87 754
rect 611 737 659 754
rect -659 642 -611 659
rect -87 642 -39 659
rect -659 611 -642 642
rect -56 611 -39 642
rect -601 105 -593 593
rect -105 105 -97 593
rect -659 56 -642 87
rect -56 56 -39 87
rect -659 39 -611 56
rect -87 39 -39 56
rect 39 642 87 659
rect 611 642 659 659
rect 39 611 56 642
rect 642 611 659 642
rect 97 105 105 593
rect 593 105 601 593
rect 39 56 56 87
rect 642 56 659 87
rect 39 39 87 56
rect 611 39 659 56
rect -659 -56 -611 -39
rect -87 -56 -39 -39
rect -659 -87 -642 -56
rect -56 -87 -39 -56
rect -601 -593 -593 -105
rect -105 -593 -97 -105
rect -659 -642 -642 -611
rect -56 -642 -39 -611
rect -659 -659 -611 -642
rect -87 -659 -39 -642
rect 39 -56 87 -39
rect 611 -56 659 -39
rect 39 -87 56 -56
rect 642 -87 659 -56
rect 97 -593 105 -105
rect 593 -593 601 -105
rect 39 -642 56 -611
rect 642 -642 659 -611
rect 39 -659 87 -642
rect 611 -659 659 -642
rect -659 -754 -611 -737
rect -87 -754 -39 -737
rect -659 -785 -642 -754
rect -56 -785 -39 -754
rect -601 -1291 -593 -803
rect -105 -1291 -97 -803
rect -659 -1340 -642 -1309
rect -56 -1340 -39 -1309
rect -659 -1357 -611 -1340
rect -87 -1357 -39 -1340
rect 39 -754 87 -737
rect 611 -754 659 -737
rect 39 -785 56 -754
rect 642 -785 659 -754
rect 97 -1291 105 -803
rect 593 -1291 601 -803
rect 39 -1340 56 -1309
rect 642 -1340 659 -1309
rect 39 -1357 87 -1340
rect 611 -1357 659 -1340
rect -659 -1452 -611 -1435
rect -87 -1452 -39 -1435
rect -659 -1483 -642 -1452
rect -56 -1483 -39 -1452
rect -601 -1989 -593 -1501
rect -105 -1989 -97 -1501
rect -659 -2038 -642 -2007
rect -56 -2038 -39 -2007
rect -659 -2055 -611 -2038
rect -87 -2055 -39 -2038
rect 39 -1452 87 -1435
rect 611 -1452 659 -1435
rect 39 -1483 56 -1452
rect 642 -1483 659 -1452
rect 97 -1989 105 -1501
rect 593 -1989 601 -1501
rect 39 -2038 56 -2007
rect 642 -2038 659 -2007
rect 39 -2055 87 -2038
rect 611 -2055 659 -2038
rect -659 -2150 -611 -2133
rect -87 -2150 -39 -2133
rect -659 -2181 -642 -2150
rect -56 -2181 -39 -2150
rect -601 -2687 -593 -2199
rect -105 -2687 -97 -2199
rect -659 -2736 -642 -2705
rect -56 -2736 -39 -2705
rect -659 -2753 -611 -2736
rect -87 -2753 -39 -2736
rect 39 -2150 87 -2133
rect 611 -2150 659 -2133
rect 39 -2181 56 -2150
rect 642 -2181 659 -2150
rect 97 -2687 105 -2199
rect 593 -2687 601 -2199
rect 39 -2736 56 -2705
rect 642 -2736 659 -2705
rect 39 -2753 87 -2736
rect 611 -2753 659 -2736
rect -764 -2841 -747 -2810
rect 747 -2841 764 -2810
rect -764 -2858 -716 -2841
rect 716 -2858 764 -2841
<< viali >>
rect -593 2199 -105 2687
rect 105 2199 593 2687
rect -593 1501 -105 1989
rect 105 1501 593 1989
rect -593 803 -105 1291
rect 105 803 593 1291
rect -593 105 -105 593
rect 105 105 593 593
rect -593 -593 -105 -105
rect 105 -593 593 -105
rect -593 -1291 -105 -803
rect 105 -1291 593 -803
rect -593 -1989 -105 -1501
rect 105 -1989 593 -1501
rect -593 -2687 -105 -2199
rect 105 -2687 593 -2199
<< metal1 >>
rect -599 2687 -99 2690
rect -599 2199 -593 2687
rect -105 2199 -99 2687
rect -599 2196 -99 2199
rect 99 2687 599 2690
rect 99 2199 105 2687
rect 593 2199 599 2687
rect 99 2196 599 2199
rect -599 1989 -99 1992
rect -599 1501 -593 1989
rect -105 1501 -99 1989
rect -599 1498 -99 1501
rect 99 1989 599 1992
rect 99 1501 105 1989
rect 593 1501 599 1989
rect 99 1498 599 1501
rect -599 1291 -99 1294
rect -599 803 -593 1291
rect -105 803 -99 1291
rect -599 800 -99 803
rect 99 1291 599 1294
rect 99 803 105 1291
rect 593 803 599 1291
rect 99 800 599 803
rect -599 593 -99 596
rect -599 105 -593 593
rect -105 105 -99 593
rect -599 102 -99 105
rect 99 593 599 596
rect 99 105 105 593
rect 593 105 599 593
rect 99 102 599 105
rect -599 -105 -99 -102
rect -599 -593 -593 -105
rect -105 -593 -99 -105
rect -599 -596 -99 -593
rect 99 -105 599 -102
rect 99 -593 105 -105
rect 593 -593 599 -105
rect 99 -596 599 -593
rect -599 -803 -99 -800
rect -599 -1291 -593 -803
rect -105 -1291 -99 -803
rect -599 -1294 -99 -1291
rect 99 -803 599 -800
rect 99 -1291 105 -803
rect 593 -1291 599 -803
rect 99 -1294 599 -1291
rect -599 -1501 -99 -1498
rect -599 -1989 -593 -1501
rect -105 -1989 -99 -1501
rect -599 -1992 -99 -1989
rect 99 -1501 599 -1498
rect 99 -1989 105 -1501
rect 593 -1989 599 -1501
rect 99 -1992 599 -1989
rect -599 -2199 -99 -2196
rect -599 -2687 -593 -2199
rect -105 -2687 -99 -2199
rect -599 -2690 -99 -2687
rect 99 -2199 599 -2196
rect 99 -2687 105 -2199
rect 593 -2687 599 -2199
rect 99 -2690 599 -2687
<< properties >>
string FIXED_BBOX 47 2141 650 2744
string gencell sky130_fd_pr__diode_pd2nw_11v0
string library sky130
string parameters w 5 l 5 area 25.0 peri 20.0 nx 2 ny 8 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 0 compatible {sky130_fd_pr__diode_pd2nw_05v5 sky130_fd_pr__diode_pd2nw_05v5_lvt  sky130_fd_pr__diode_pd2nw_05v5_hvt sky130_fd_pr__diode_pd2nw_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
