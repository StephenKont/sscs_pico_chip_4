magic
tech sky130A
timestamp 1665661446
<< metal3 >>
rect -575 -550 524 550
<< mimcap >>
rect -525 480 475 500
rect -525 -480 -505 480
rect 455 -480 475 480
rect -525 -500 475 -480
<< mimcapcontact >>
rect -505 -480 455 480
<< properties >>
string FIXED_BBOX -575 -550 525 550
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10 l 10 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
