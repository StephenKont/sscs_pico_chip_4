magic
tech sky130A
timestamp 1666550119
<< metal4 >>
rect -1541 3650 -1371 3692
rect 1115 3650 1285 3674
rect -2656 2819 -158 3650
rect 5 2819 2502 3650
rect -2656 2545 2502 2819
rect -2656 1250 -158 2545
rect 5 1250 2502 2545
rect -1541 1200 -1371 1250
rect 1115 1200 1285 1250
rect -2656 53 -159 1200
rect 5 53 2502 1200
rect -2656 -221 2502 53
rect -2656 -1200 -159 -221
rect 5 -1200 2502 -221
rect -1541 -1250 -1371 -1200
rect 1115 -1250 1285 -1200
rect -2656 -2282 -161 -1250
rect 6 -2282 2502 -1250
rect -2656 -2556 2502 -2282
rect -2656 -3650 -161 -2556
rect 6 -3650 2502 -2556
rect -1541 -3664 -1371 -3650
rect 1115 -3682 1285 -3650
<< mimcap2 >>
rect -2606 3580 -306 3600
rect -2606 1320 -2586 3580
rect -326 1320 -306 3580
rect -2606 1300 -306 1320
rect 55 3580 2355 3600
rect 55 1320 75 3580
rect 2335 1320 2355 3580
rect 55 1300 2355 1320
rect -2606 1130 -306 1150
rect -2606 -1130 -2586 1130
rect -326 -1130 -306 1130
rect -2606 -1150 -306 -1130
rect 55 1130 2355 1150
rect 55 -1130 75 1130
rect 2335 -1130 2355 1130
rect 55 -1150 2355 -1130
rect -2606 -1320 -306 -1300
rect -2606 -3580 -2586 -1320
rect -326 -3580 -306 -1320
rect -2606 -3600 -306 -3580
rect 55 -1320 2355 -1300
rect 55 -3580 75 -1320
rect 2335 -3580 2355 -1320
rect 55 -3600 2355 -3580
<< mimcap2contact >>
rect -2586 1320 -326 3580
rect 75 1320 2335 3580
rect -2586 -1130 -326 1130
rect 75 -1130 2335 1130
rect -2586 -3580 -326 -1320
rect 75 -3580 2335 -1320
<< metal5 >>
rect -1536 3592 -1376 3675
rect -326 3592 -166 3675
rect 1125 3592 1285 3675
rect 2335 3592 2495 3675
rect -2598 3580 -166 3592
rect -2598 1320 -2586 3580
rect -326 2817 -166 3580
rect 63 3580 2495 3592
rect 63 2817 75 3580
rect -326 2544 75 2817
rect -326 1320 -166 2544
rect -2598 1308 -166 1320
rect 63 1320 75 2544
rect 2335 1320 2495 3580
rect 63 1308 2495 1320
rect -1536 1142 -1376 1308
rect -326 1142 -166 1308
rect 1125 1142 1285 1308
rect 2335 1142 2495 1308
rect -2598 1130 -166 1142
rect -2598 -1130 -2586 1130
rect -326 49 -166 1130
rect 63 1130 2495 1142
rect 63 49 75 1130
rect -326 -224 75 49
rect -326 -1130 -166 -224
rect -2598 -1142 -166 -1130
rect 63 -1130 75 -224
rect 2335 -1130 2495 1130
rect 63 -1142 2495 -1130
rect -1536 -1308 -1376 -1142
rect -326 -1308 -166 -1142
rect 1125 -1308 1285 -1142
rect 2335 -1308 2495 -1142
rect -2598 -1320 -166 -1308
rect -2598 -3580 -2586 -1320
rect -326 -2280 -166 -1320
rect 63 -1320 2495 -1308
rect 63 -2280 75 -1320
rect -326 -2553 75 -2280
rect -326 -3580 -166 -2553
rect -2598 -3592 -166 -3580
rect 63 -3580 75 -2553
rect 2335 -3580 2495 -1320
rect 63 -3592 2495 -3580
rect -1536 -3675 -1376 -3592
rect -326 -3675 -166 -3592
rect 1125 -3675 1285 -3592
rect 2335 -3675 2495 -3592
<< properties >>
string FIXED_BBOX 5 1250 2405 3650
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 23.00 l 23.00 val 1.075k carea 2.00 cperi 0.19 nx 2 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
