magic
tech sky130A
magscale 1 2
timestamp 1669392366
<< locali >>
rect 556599 154474 556632 154508
rect 556599 153142 556632 153176
rect 53408 130140 53902 130170
rect 53408 128994 53436 130140
rect 53868 128994 53902 130140
rect 53408 128970 53902 128994
rect 62794 127656 63358 127692
rect 62794 126510 62876 127656
rect 63308 126510 63358 127656
rect 62794 126478 63358 126510
rect 53408 126178 53902 126208
rect 53408 125032 53436 126178
rect 53868 125032 53902 126178
rect 53408 125008 53902 125032
rect 62794 123694 63358 123730
rect 62794 122548 62876 123694
rect 63308 122548 63358 123694
rect 62794 122516 63358 122548
rect 53408 122216 53902 122246
rect 53408 121070 53436 122216
rect 53868 121070 53902 122216
rect 53408 121046 53902 121070
rect 62794 119732 63358 119768
rect 62794 118586 62876 119732
rect 63308 118586 63358 119732
rect 62794 118554 63358 118586
rect 53408 118254 53902 118284
rect 53408 117108 53436 118254
rect 53868 117108 53902 118254
rect 53408 117084 53902 117108
rect 62794 115770 63358 115806
rect 62794 114624 62876 115770
rect 63308 114624 63358 115770
rect 62794 114592 63358 114624
<< viali >>
rect 467844 450395 468039 450429
rect 468206 450395 468402 450429
rect 468844 450395 469039 450429
rect 469206 450395 469402 450429
rect 467748 449775 467782 450333
rect 468054 450185 468192 450219
rect 467958 449985 467992 450123
rect 468090 450021 468156 450087
rect 468254 449985 468288 450123
rect 468464 449775 468498 450333
rect 468748 449775 468782 450333
rect 469054 450185 469192 450219
rect 468958 449985 468992 450123
rect 469090 450021 469156 450087
rect 469254 449985 469288 450123
rect 469464 449775 469498 450333
rect 467844 449679 468402 449713
rect 468844 449679 469402 449713
rect 334420 389741 334615 389775
rect 334782 389741 334978 389775
rect 335420 389741 335615 389775
rect 335782 389741 335978 389775
rect 334324 389121 334358 389679
rect 334630 389531 334768 389565
rect 334534 389331 334568 389469
rect 334830 389331 334864 389469
rect 335040 389121 335074 389679
rect 335324 389121 335358 389679
rect 335630 389531 335768 389565
rect 335534 389331 335568 389469
rect 335830 389331 335864 389469
rect 336040 389121 336074 389679
rect 334420 389025 334978 389059
rect 335420 389025 335978 389059
rect 554342 154476 555336 154510
rect 555946 154474 556599 154508
rect 553707 154337 554081 154371
rect 553611 153897 553645 154275
rect 554143 153897 554177 154275
rect 553707 153801 554081 153835
rect 553707 153695 554081 153729
rect 553611 153255 553645 153633
rect 554143 153255 554177 153633
rect 554246 153240 554280 154414
rect 555398 153240 555432 154414
rect 555850 153238 555884 154412
rect 556654 153238 556688 154412
rect 553707 153159 554081 153193
rect 554342 153144 555336 153178
rect 555946 153142 556599 153176
rect 554208 152874 555510 152908
rect 556186 152874 556448 152908
rect 553694 152808 553950 152842
rect 553598 152368 553632 152746
rect 554012 152368 554046 152746
rect 553694 152272 553950 152306
rect 553694 152166 553950 152200
rect 553598 151726 553632 152104
rect 554012 151726 554046 152104
rect 553694 151630 553950 151664
rect 554112 151656 554146 152812
rect 555572 151656 555606 152812
rect 556090 151656 556124 152812
rect 556510 151656 556544 152812
rect 554208 151560 555510 151594
rect 556186 151560 556448 151594
rect 57842 148102 58098 148136
rect 58362 148102 58618 148136
rect 58882 148102 59138 148136
rect 59402 148102 59658 148136
rect 57746 147312 57780 148040
rect 58160 147312 58194 148040
rect 58266 147312 58300 148040
rect 58680 147312 58714 148040
rect 58786 147312 58820 148040
rect 59200 147312 59234 148040
rect 59306 147312 59340 148040
rect 59720 147312 59754 148040
rect 57842 147216 58098 147250
rect 58362 147216 58618 147250
rect 58882 147216 59138 147250
rect 59402 147216 59658 147250
rect 551479 147089 551674 147123
rect 551841 147089 552037 147123
rect 552479 147089 552674 147123
rect 552841 147089 553037 147123
rect 551383 146469 551417 147027
rect 551689 146879 551827 146913
rect 551593 146679 551627 146817
rect 551725 146715 551791 146781
rect 551889 146679 551923 146817
rect 552099 146469 552133 147027
rect 552383 146469 552417 147027
rect 552689 146879 552827 146913
rect 552593 146679 552627 146817
rect 552725 146715 552791 146781
rect 552889 146679 552923 146817
rect 553099 146469 553133 147027
rect 551479 146373 552037 146407
rect 552479 146373 553037 146407
rect 60480 146119 60675 146153
rect 60842 146119 61038 146153
rect 61480 146119 61675 146153
rect 61842 146119 62038 146153
rect 62480 146119 62675 146153
rect 62842 146119 63038 146153
rect 63480 146119 63675 146153
rect 63842 146119 64038 146153
rect 53732 146030 53927 146064
rect 54094 146030 54290 146064
rect 54732 146030 54927 146064
rect 55094 146030 55290 146064
rect 55732 146030 55927 146064
rect 56094 146030 56290 146064
rect 56732 146030 56927 146064
rect 57094 146030 57290 146064
rect 53636 145410 53670 145968
rect 53942 145820 54080 145854
rect 53846 145620 53880 145758
rect 53978 145656 54044 145722
rect 54142 145620 54176 145758
rect 54352 145410 54386 145968
rect 54636 145410 54670 145968
rect 54942 145820 55080 145854
rect 54846 145620 54880 145758
rect 54978 145656 55044 145722
rect 55142 145620 55176 145758
rect 55352 145410 55386 145968
rect 55636 145410 55670 145968
rect 55942 145820 56080 145854
rect 55846 145620 55880 145758
rect 55978 145656 56044 145722
rect 56142 145620 56176 145758
rect 56352 145410 56386 145968
rect 56636 145410 56670 145968
rect 56942 145820 57080 145854
rect 56846 145620 56880 145758
rect 56978 145656 57044 145722
rect 57142 145620 57176 145758
rect 57352 145410 57386 145968
rect 60384 145499 60418 146057
rect 60690 145909 60828 145943
rect 60594 145709 60628 145847
rect 60726 145745 60792 145811
rect 60890 145709 60924 145847
rect 61100 145499 61134 146057
rect 61384 145499 61418 146057
rect 61690 145909 61828 145943
rect 61594 145709 61628 145847
rect 61726 145745 61792 145811
rect 61890 145709 61924 145847
rect 62100 145499 62134 146057
rect 62384 145499 62418 146057
rect 62690 145909 62828 145943
rect 62594 145709 62628 145847
rect 62726 145745 62792 145811
rect 62890 145709 62924 145847
rect 63100 145499 63134 146057
rect 63384 145499 63418 146057
rect 63690 145909 63828 145943
rect 63594 145709 63628 145847
rect 63726 145745 63792 145811
rect 63890 145709 63924 145847
rect 64100 145499 64134 146057
rect 60480 145403 61038 145437
rect 61480 145403 62038 145437
rect 62480 145403 63038 145437
rect 63480 145403 64038 145437
rect 53732 145314 54290 145348
rect 54732 145314 55290 145348
rect 55732 145314 56290 145348
rect 56732 145314 57290 145348
rect 53402 130236 63342 130270
rect 53306 126476 53340 130174
rect 53436 128994 53868 130140
rect 62876 126510 63308 127656
rect 63404 126476 63438 130174
rect 53402 126380 63342 126414
rect 53402 126274 63342 126308
rect 53306 122514 53340 126212
rect 53436 125032 53868 126178
rect 62876 122548 63308 123694
rect 63404 122514 63438 126212
rect 53402 122418 63342 122452
rect 53402 122312 63342 122346
rect 53306 118552 53340 122250
rect 53436 121070 53868 122216
rect 62876 118586 63308 119732
rect 63404 118552 63438 122250
rect 53402 118456 63342 118490
rect 53402 118350 63342 118384
rect 53306 114590 53340 118288
rect 53436 117108 53868 118254
rect 62876 114624 63308 115770
rect 63404 114590 63438 118288
rect 53402 114494 63342 114528
<< metal1 >>
rect 351259 697923 404827 699695
rect 406599 697923 406605 699695
rect 145394 681965 165394 682901
rect 145394 674731 146520 681965
rect 164088 674731 165394 681965
rect 145394 567969 165394 674731
rect 351259 610221 353031 697923
rect 529662 696917 530093 696928
rect 529662 696526 529691 696917
rect 530082 696526 533502 696917
rect 529662 696509 530093 696526
rect 418923 692927 531009 693157
rect 418923 690516 419153 692927
rect 418001 690286 419153 690516
rect 530779 685003 531009 692927
rect 533111 691809 533502 696526
rect 533111 691418 535568 691809
rect 540110 687288 540426 687322
rect 540110 687119 540137 687288
rect 540399 687119 540426 687288
rect 540110 687092 540426 687119
rect 540143 685003 540373 687092
rect 530779 684773 540373 685003
rect 540143 684600 540373 684773
rect 540143 684370 579810 684600
rect 442918 679662 462918 680730
rect 442918 669616 443952 679662
rect 462134 669616 462918 679662
rect 442918 613648 462918 669616
rect 442918 599950 444062 613648
rect 461834 599950 462918 613648
rect 442918 598730 462918 599950
rect 579580 583727 579810 684370
rect 579559 583706 579826 583727
rect 579559 583476 579580 583706
rect 579810 583476 579826 583706
rect 579559 583451 579826 583476
rect 145394 556095 146784 567969
rect 164076 556095 165394 567969
rect 145394 553901 165394 556095
rect 145398 511617 165398 512901
rect 145398 498073 146694 511617
rect 163458 498073 165398 511617
rect 145398 409147 165398 498073
rect 468092 460164 468156 460170
rect 467736 450441 468045 450442
rect 467735 450429 468045 450441
rect 467735 450395 467844 450429
rect 468039 450395 468045 450429
rect 467735 450383 468045 450395
rect 467735 450333 467794 450383
rect 467735 449775 467748 450333
rect 467782 449775 467794 450333
rect 468092 450231 468156 460100
rect 469092 458678 469156 458684
rect 468200 450429 468510 450442
rect 468736 450441 469045 450442
rect 468200 450395 468206 450429
rect 468402 450395 468510 450429
rect 468200 450383 468510 450395
rect 468452 450333 468510 450383
rect 467946 450219 468300 450231
rect 467946 450185 468054 450219
rect 468192 450185 468300 450219
rect 467946 450173 468300 450185
rect 467946 450123 468004 450173
rect 467946 449985 467958 450123
rect 467992 449985 468004 450123
rect 468242 450123 468300 450173
rect 467946 449877 468004 449985
rect 468078 450087 468168 450099
rect 468078 450021 468090 450087
rect 468156 450021 468168 450087
rect 467735 449725 467794 449775
rect 468078 449725 468168 450021
rect 468242 449985 468254 450123
rect 468288 449985 468300 450123
rect 468242 449877 468300 449985
rect 468452 449775 468464 450333
rect 468498 449775 468510 450333
rect 468452 449725 468510 449775
rect 467735 449713 468510 449725
rect 467735 449679 467844 449713
rect 468402 449679 468510 449713
rect 467735 449667 468510 449679
rect 467735 449521 467794 449667
rect 468452 449521 468510 449667
rect 468735 450429 469045 450441
rect 468735 450395 468844 450429
rect 469039 450395 469045 450429
rect 468735 450383 469045 450395
rect 468735 450333 468794 450383
rect 468735 449775 468748 450333
rect 468782 449775 468794 450333
rect 469092 450231 469156 458614
rect 469200 450429 469510 450442
rect 469200 450395 469206 450429
rect 469402 450395 469510 450429
rect 469200 450383 469510 450395
rect 469452 450333 469510 450383
rect 468946 450219 469300 450231
rect 468946 450185 469054 450219
rect 469192 450185 469300 450219
rect 468946 450173 469300 450185
rect 468946 450123 469004 450173
rect 468946 449985 468958 450123
rect 468992 449985 469004 450123
rect 469242 450123 469300 450173
rect 468946 449877 469004 449985
rect 469078 450087 469168 450099
rect 469078 450021 469090 450087
rect 469156 450021 469168 450087
rect 468735 449725 468794 449775
rect 469078 449725 469168 450021
rect 469242 449985 469254 450123
rect 469288 449985 469300 450123
rect 469242 449877 469300 449985
rect 469452 449775 469464 450333
rect 469498 449775 469510 450333
rect 469452 449725 469510 449775
rect 468735 449713 469510 449725
rect 468735 449679 468844 449713
rect 469402 449679 469510 449713
rect 468735 449667 469510 449679
rect 468735 449521 468794 449667
rect 469452 449521 469510 449667
rect 467580 449507 469674 449521
rect 467580 449422 467592 449507
rect 469659 449422 469674 449507
rect 467580 449411 469674 449422
rect 145398 401839 146500 409147
rect 164068 401839 165398 409147
rect 145398 400903 165398 401839
rect 335657 390802 335741 390811
rect 335657 390738 335668 390802
rect 335732 390738 335741 390802
rect 335657 390728 335741 390738
rect 334650 390146 334758 390164
rect 334650 390082 334668 390146
rect 334732 390082 334758 390146
rect 334650 390066 334758 390082
rect 334312 389787 334621 389788
rect 334311 389775 334621 389787
rect 334311 389741 334420 389775
rect 334615 389741 334621 389775
rect 334311 389729 334621 389741
rect 334311 389679 334370 389729
rect 334311 389121 334324 389679
rect 334358 389121 334370 389679
rect 334668 389577 334732 390066
rect 334776 389775 335086 389788
rect 335312 389787 335621 389788
rect 334776 389741 334782 389775
rect 334978 389741 335086 389775
rect 334776 389729 335086 389741
rect 335028 389679 335086 389729
rect 334522 389565 334876 389577
rect 334522 389531 334630 389565
rect 334768 389531 334876 389565
rect 334522 389519 334876 389531
rect 334522 389469 334580 389519
rect 334522 389331 334534 389469
rect 334568 389331 334580 389469
rect 334818 389469 334876 389519
rect 334522 389223 334580 389331
rect 334311 389071 334370 389121
rect 334654 389071 334744 389445
rect 334818 389331 334830 389469
rect 334864 389331 334876 389469
rect 334818 389223 334876 389331
rect 335028 389121 335040 389679
rect 335074 389121 335086 389679
rect 335028 389071 335086 389121
rect 334311 389059 335086 389071
rect 334311 389025 334420 389059
rect 334978 389025 335086 389059
rect 334311 389013 335086 389025
rect 334311 388853 334370 389013
rect 335028 388853 335086 389013
rect 335311 389775 335621 389787
rect 335311 389741 335420 389775
rect 335615 389741 335621 389775
rect 335311 389729 335621 389741
rect 335311 389679 335370 389729
rect 335311 389121 335324 389679
rect 335358 389121 335370 389679
rect 335668 389577 335732 390728
rect 335776 389775 336086 389788
rect 335776 389741 335782 389775
rect 335978 389741 336086 389775
rect 335776 389729 336086 389741
rect 336028 389679 336086 389729
rect 335522 389565 335876 389577
rect 335522 389531 335630 389565
rect 335768 389531 335876 389565
rect 335522 389519 335876 389531
rect 335522 389469 335580 389519
rect 335522 389331 335534 389469
rect 335568 389331 335580 389469
rect 335818 389469 335876 389519
rect 335522 389223 335580 389331
rect 335311 389071 335370 389121
rect 335654 389071 335744 389445
rect 335818 389331 335830 389469
rect 335864 389331 335876 389469
rect 335818 389223 335876 389331
rect 336028 389121 336040 389679
rect 336074 389121 336086 389679
rect 336028 389071 336086 389121
rect 335311 389059 336086 389071
rect 335311 389025 335420 389059
rect 335978 389025 336086 389059
rect 335311 389013 336086 389025
rect 335311 388853 335370 389013
rect 336028 388853 336086 389013
rect 333727 388772 336528 388853
rect 333727 387884 333824 388772
rect 336416 387884 336528 388772
rect 333727 387811 336528 387884
rect 550243 155139 550317 155145
rect 550317 155065 554813 155139
rect 550243 155059 550317 155065
rect 554739 154546 554813 155065
rect 554210 154510 556724 154546
rect 554210 154482 554342 154510
rect 554208 154476 554342 154482
rect 555336 154508 556724 154510
rect 555336 154476 555946 154508
rect 554208 154474 555946 154476
rect 556599 154474 556724 154508
rect 554208 154460 556724 154474
rect 554208 154414 554298 154460
rect 554208 154408 554246 154414
rect 553574 154371 554246 154408
rect 553574 154337 553707 154371
rect 554081 154337 554246 154371
rect 553574 154322 554246 154337
rect 553574 154275 553660 154322
rect 553574 153897 553611 154275
rect 553645 153897 553660 154275
rect 553794 154275 553994 154282
rect 553794 154223 553806 154275
rect 553982 154223 553994 154275
rect 553794 154217 553994 154223
rect 554128 154275 554246 154322
rect 553707 154195 553771 154201
rect 553707 153977 553713 154195
rect 553765 153977 553771 154195
rect 553707 153971 553771 153977
rect 553574 153850 553660 153897
rect 553804 153949 554004 153956
rect 553804 153897 553816 153949
rect 553992 153897 554004 153949
rect 553804 153891 554004 153897
rect 554128 153897 554143 154275
rect 554177 153897 554246 154275
rect 554128 153850 554246 153897
rect 553574 153835 554246 153850
rect 553574 153801 553707 153835
rect 554081 153801 554246 153835
rect 553574 153729 554246 153801
rect 553574 153695 553707 153729
rect 554081 153695 554246 153729
rect 553574 153680 554246 153695
rect 553574 153633 553660 153680
rect 553574 153255 553611 153633
rect 553645 153255 553660 153633
rect 553804 153633 554004 153640
rect 553804 153581 553817 153633
rect 553993 153581 554004 153633
rect 553804 153575 554004 153581
rect 554128 153633 554246 153680
rect 553707 153553 553771 153559
rect 553707 153335 553713 153553
rect 553765 153335 553771 153553
rect 553707 153329 553771 153335
rect 553574 153208 553660 153255
rect 553803 153307 554003 153313
rect 553803 153255 553815 153307
rect 553991 153255 554003 153307
rect 553803 153248 554003 153255
rect 554128 153255 554143 153633
rect 554177 153255 554246 153633
rect 554128 153240 554246 153255
rect 554280 153240 554298 154414
rect 555378 154414 555468 154460
rect 554348 154316 554411 154327
rect 554348 153333 554354 154316
rect 554406 153333 554411 154316
rect 554961 154316 555024 154327
rect 554348 153327 554411 153333
rect 554650 153581 554721 153590
rect 554650 153337 554659 153581
rect 554711 153337 554721 153581
rect 554650 153327 554721 153337
rect 554961 153333 554967 154316
rect 555019 153333 555024 154316
rect 554961 153327 555024 153333
rect 555259 153578 555335 153590
rect 555259 153334 555269 153578
rect 555325 153334 555335 153578
rect 555259 153325 555335 153334
rect 554128 153208 554298 153240
rect 554404 153288 555272 153294
rect 554404 153236 554410 153288
rect 555264 153236 555272 153288
rect 554404 153230 555272 153236
rect 555378 153240 555398 154414
rect 555432 153240 555468 154414
rect 553574 153193 554298 153208
rect 553574 153159 553707 153193
rect 554081 153192 554298 153193
rect 555378 153192 555468 153240
rect 555814 154412 555904 154460
rect 555814 153238 555850 154412
rect 555884 153238 555904 154412
rect 556086 154425 556542 154431
rect 556086 154372 556092 154425
rect 556536 154372 556542 154425
rect 556086 154366 556542 154372
rect 556634 154412 556724 154460
rect 555948 154318 556010 154325
rect 555948 153331 555954 154318
rect 556006 153331 556010 154318
rect 555948 153325 556010 153331
rect 556044 154318 556106 154325
rect 556044 153331 556050 154318
rect 556102 153331 556106 154318
rect 556044 153325 556106 153331
rect 556140 154318 556202 154325
rect 556140 153331 556146 154318
rect 556198 153331 556202 154318
rect 556140 153325 556202 153331
rect 556236 154318 556298 154325
rect 556236 153331 556242 154318
rect 556294 153331 556298 154318
rect 556236 153325 556298 153331
rect 556332 154318 556394 154325
rect 556332 153331 556338 154318
rect 556390 153331 556394 154318
rect 556332 153325 556394 153331
rect 556428 154318 556490 154325
rect 556428 153331 556434 154318
rect 556486 153331 556490 154318
rect 556428 153325 556490 153331
rect 556524 154318 556586 154325
rect 556524 153331 556530 154318
rect 556582 153331 556586 154318
rect 556524 153325 556586 153331
rect 555814 153192 555904 153238
rect 555996 153278 556446 153284
rect 555996 153226 556019 153278
rect 556436 153226 556446 153278
rect 555996 153220 556446 153226
rect 556634 153238 556654 154412
rect 556688 153238 556724 154412
rect 556634 153192 556724 153238
rect 554081 153178 556724 153192
rect 554081 153159 554342 153178
rect 553574 153144 554342 153159
rect 555336 153176 556724 153178
rect 555336 153144 555946 153176
rect 553574 153142 555946 153144
rect 556599 153142 556724 153176
rect 553574 153122 556724 153142
rect 554208 153106 556724 153122
rect 554076 152908 556580 152944
rect 554076 152878 554208 152908
rect 553562 152874 554208 152878
rect 555510 152874 556186 152908
rect 556448 152874 556580 152908
rect 553562 152860 556580 152874
rect 553562 152842 554160 152860
rect 553562 152808 553694 152842
rect 553950 152812 554160 152842
rect 555558 152858 556580 152860
rect 553950 152808 554112 152812
rect 553562 152794 554112 152808
rect 553562 152746 553648 152794
rect 553562 152368 553598 152746
rect 553632 152368 553648 152746
rect 553779 152746 553875 152756
rect 553779 152694 553786 152746
rect 553867 152694 553875 152746
rect 553779 152688 553875 152694
rect 553996 152746 554112 152794
rect 553684 152666 553748 152673
rect 553684 152448 553690 152666
rect 553742 152448 553748 152666
rect 553684 152442 553748 152448
rect 553562 152322 553648 152368
rect 553779 152419 553875 152426
rect 553779 152367 553787 152419
rect 553868 152367 553875 152419
rect 553779 152358 553875 152367
rect 553996 152368 554012 152746
rect 554046 152368 554112 152746
rect 553996 152322 554112 152368
rect 553562 152306 554112 152322
rect 553562 152272 553694 152306
rect 553950 152272 554112 152306
rect 553562 152200 554112 152272
rect 553562 152166 553694 152200
rect 553950 152166 554112 152200
rect 553562 152146 554112 152166
rect 553562 152104 553648 152146
rect 553562 151726 553598 152104
rect 553632 151726 553648 152104
rect 553780 152105 553876 152114
rect 553780 152053 553788 152105
rect 553869 152053 553876 152105
rect 553780 152046 553876 152053
rect 553996 152104 554112 152146
rect 553684 152024 553748 152030
rect 553684 151806 553690 152024
rect 553742 151806 553748 152024
rect 553684 151799 553748 151806
rect 553562 151680 553648 151726
rect 553780 151777 553876 151785
rect 553780 151725 553787 151777
rect 553868 151725 553876 151777
rect 553780 151717 553876 151725
rect 553996 151726 554012 152104
rect 554046 151726 554112 152104
rect 553996 151680 554112 151726
rect 553562 151664 554112 151680
rect 553562 151630 553694 151664
rect 553950 151656 554112 151664
rect 554146 151656 554160 152812
rect 554272 152820 555446 152826
rect 554272 152768 554277 152820
rect 555439 152768 555446 152820
rect 554272 152762 555446 152768
rect 555558 152812 555642 152858
rect 554214 152722 554282 152734
rect 554214 151746 554226 152722
rect 554278 151746 554282 152722
rect 554502 152728 554593 152734
rect 554502 152349 554520 152728
rect 554583 152349 554593 152728
rect 554502 152329 554593 152349
rect 554824 152717 554892 152734
rect 554214 151734 554282 151746
rect 554824 151741 554834 152717
rect 554886 151741 554892 152717
rect 555119 152727 555216 152734
rect 555119 152348 555135 152727
rect 555198 152348 555216 152727
rect 555119 152325 555216 152348
rect 555438 152717 555506 152734
rect 554824 151734 554892 151741
rect 555438 151741 555446 152717
rect 555498 151741 555506 152717
rect 555438 151734 555506 151741
rect 553950 151630 554160 151656
rect 553562 151608 554160 151630
rect 555558 151656 555572 152812
rect 555606 151656 555642 152812
rect 555558 151608 555642 151656
rect 556054 152812 556138 152858
rect 556054 151656 556090 152812
rect 556124 151656 556138 152812
rect 556250 152824 556432 152830
rect 556250 152772 556266 152824
rect 556416 152772 556432 152824
rect 556250 152766 556432 152772
rect 556496 152812 556580 152858
rect 556192 152727 556255 152734
rect 556192 151742 556197 152727
rect 556249 151742 556255 152727
rect 556192 151734 556255 151742
rect 556289 152727 556350 152734
rect 556289 151740 556293 152727
rect 556345 151740 556350 152727
rect 556289 151734 556350 151740
rect 556392 152727 556454 152734
rect 556392 151742 556397 152727
rect 556449 151742 556454 152727
rect 556392 151734 556454 151742
rect 556054 151608 556138 151656
rect 556216 151696 556302 151702
rect 556216 151644 556223 151696
rect 556294 151644 556302 151696
rect 556216 151638 556302 151644
rect 556496 151656 556510 152812
rect 556544 151656 556580 152812
rect 556496 151608 556580 151656
rect 553562 151594 556580 151608
rect 554076 151560 554208 151594
rect 555510 151560 556186 151594
rect 556448 151560 556580 151594
rect 554076 151524 556580 151560
rect 59223 150309 59229 150383
rect 59303 150309 60774 150383
rect 554693 150383 554767 151524
rect 61274 150309 554767 150383
rect 53980 148852 59506 148916
rect 59570 148852 59576 148916
rect 53624 146076 53933 146077
rect 53623 146064 53933 146076
rect 53623 146030 53732 146064
rect 53927 146030 53933 146064
rect 53623 146018 53933 146030
rect 53623 145968 53682 146018
rect 53623 145410 53636 145968
rect 53670 145410 53682 145968
rect 53980 145866 54044 148852
rect 54980 148640 58986 148704
rect 59050 148640 59056 148704
rect 59638 148682 59644 148746
rect 59708 148682 63792 148746
rect 54088 146064 54398 146077
rect 54624 146076 54933 146077
rect 54088 146030 54094 146064
rect 54290 146030 54398 146064
rect 54088 146018 54398 146030
rect 54340 145968 54398 146018
rect 53834 145854 54188 145866
rect 53834 145820 53942 145854
rect 54080 145820 54188 145854
rect 53834 145808 54188 145820
rect 53834 145758 53892 145808
rect 53834 145620 53846 145758
rect 53880 145620 53892 145758
rect 54130 145758 54188 145808
rect 53834 145512 53892 145620
rect 53966 145722 54056 145734
rect 53966 145656 53978 145722
rect 54044 145656 54056 145722
rect 53623 145360 53682 145410
rect 53966 145360 54056 145656
rect 54130 145620 54142 145758
rect 54176 145620 54188 145758
rect 54130 145512 54188 145620
rect 54340 145410 54352 145968
rect 54386 145410 54398 145968
rect 54340 145360 54398 145410
rect 53623 145348 54398 145360
rect 53623 145314 53732 145348
rect 54290 145314 54398 145348
rect 53623 145302 54398 145314
rect 53623 145219 53682 145302
rect 54340 145219 54398 145302
rect 54623 146064 54933 146076
rect 54623 146030 54732 146064
rect 54927 146030 54933 146064
rect 54623 146018 54933 146030
rect 54623 145968 54682 146018
rect 54623 145410 54636 145968
rect 54670 145410 54682 145968
rect 54980 145866 55044 148640
rect 59114 148616 59178 148622
rect 59178 148552 62792 148616
rect 59114 148546 59178 148552
rect 55980 148464 58462 148528
rect 58526 148464 58532 148528
rect 55088 146064 55398 146077
rect 55624 146076 55933 146077
rect 55088 146030 55094 146064
rect 55290 146030 55398 146064
rect 55088 146018 55398 146030
rect 55340 145968 55398 146018
rect 54834 145854 55188 145866
rect 54834 145820 54942 145854
rect 55080 145820 55188 145854
rect 54834 145808 55188 145820
rect 54834 145758 54892 145808
rect 54834 145620 54846 145758
rect 54880 145620 54892 145758
rect 55130 145758 55188 145808
rect 54834 145512 54892 145620
rect 54966 145722 55056 145734
rect 54966 145656 54978 145722
rect 55044 145656 55056 145722
rect 54623 145360 54682 145410
rect 54966 145360 55056 145656
rect 55130 145620 55142 145758
rect 55176 145620 55188 145758
rect 55130 145512 55188 145620
rect 55340 145410 55352 145968
rect 55386 145410 55398 145968
rect 55340 145360 55398 145410
rect 54623 145348 55398 145360
rect 54623 145314 54732 145348
rect 55290 145314 55398 145348
rect 54623 145302 55398 145314
rect 54623 145219 54682 145302
rect 55340 145219 55398 145302
rect 55623 146064 55933 146076
rect 55623 146030 55732 146064
rect 55927 146030 55933 146064
rect 55623 146018 55933 146030
rect 55623 145968 55682 146018
rect 55623 145410 55636 145968
rect 55670 145410 55682 145968
rect 55980 145866 56044 148464
rect 58584 148418 58590 148482
rect 58654 148418 61792 148482
rect 56980 148292 57942 148356
rect 58006 148292 58012 148356
rect 56088 146064 56398 146077
rect 56624 146076 56933 146077
rect 56088 146030 56094 146064
rect 56290 146030 56398 146064
rect 56088 146018 56398 146030
rect 56340 145968 56398 146018
rect 55834 145854 56188 145866
rect 55834 145820 55942 145854
rect 56080 145820 56188 145854
rect 55834 145808 56188 145820
rect 55834 145758 55892 145808
rect 55834 145620 55846 145758
rect 55880 145620 55892 145758
rect 56130 145758 56188 145808
rect 55834 145512 55892 145620
rect 55966 145722 56056 145734
rect 55966 145656 55978 145722
rect 56044 145656 56056 145722
rect 55623 145360 55682 145410
rect 55966 145360 56056 145656
rect 56130 145620 56142 145758
rect 56176 145620 56188 145758
rect 56130 145512 56188 145620
rect 56340 145410 56352 145968
rect 56386 145410 56398 145968
rect 56340 145360 56398 145410
rect 55623 145348 56398 145360
rect 55623 145314 55732 145348
rect 56290 145314 56398 145348
rect 55623 145302 56398 145314
rect 55623 145219 55682 145302
rect 56340 145219 56398 145302
rect 56623 146064 56933 146076
rect 56623 146030 56732 146064
rect 56927 146030 56933 146064
rect 56623 146018 56933 146030
rect 56623 145968 56682 146018
rect 56623 145410 56636 145968
rect 56670 145410 56682 145968
rect 56980 145866 57044 148292
rect 58072 148222 58078 148286
rect 58142 148222 60792 148286
rect 57710 148144 59790 148172
rect 57708 148136 59790 148144
rect 57708 148102 57842 148136
rect 58098 148102 58362 148136
rect 58618 148102 58882 148136
rect 59138 148102 59402 148136
rect 59658 148102 59790 148136
rect 57708 148092 59790 148102
rect 57708 148040 57790 148092
rect 57708 147312 57746 148040
rect 57780 147312 57790 148040
rect 57920 148042 58020 148050
rect 57920 147988 57928 148042
rect 58010 147988 58020 148042
rect 57920 147982 58020 147988
rect 58148 148040 58312 148092
rect 58052 147968 58116 147976
rect 58052 147392 58058 147968
rect 58110 147392 58116 147968
rect 58052 147376 58116 147392
rect 57708 147260 57790 147312
rect 57920 147260 58020 147370
rect 58148 147312 58160 148040
rect 58194 147312 58266 148040
rect 58300 147312 58312 148040
rect 58440 148042 58540 148050
rect 58440 147988 58448 148042
rect 58530 147988 58540 148042
rect 58440 147982 58540 147988
rect 58668 148040 58832 148092
rect 58572 147968 58636 147976
rect 58572 147392 58578 147968
rect 58630 147392 58636 147968
rect 58572 147376 58636 147392
rect 58148 147260 58312 147312
rect 58440 147260 58540 147370
rect 58668 147312 58680 148040
rect 58714 147312 58786 148040
rect 58820 147312 58832 148040
rect 58960 148042 59060 148050
rect 58960 147988 58968 148042
rect 59050 147988 59060 148042
rect 58960 147982 59060 147988
rect 59188 148040 59352 148092
rect 59092 147968 59156 147976
rect 59092 147392 59098 147968
rect 59150 147392 59156 147968
rect 59092 147376 59156 147392
rect 58668 147260 58832 147312
rect 58960 147260 59060 147370
rect 59188 147312 59200 148040
rect 59234 147312 59306 148040
rect 59340 147312 59352 148040
rect 59480 148042 59580 148050
rect 59480 147988 59488 148042
rect 59570 147988 59580 148042
rect 59480 147982 59580 147988
rect 59708 148040 59790 148092
rect 59612 147968 59676 147976
rect 59612 147392 59618 147968
rect 59670 147392 59676 147968
rect 59612 147376 59676 147392
rect 59188 147260 59352 147312
rect 59480 147260 59580 147370
rect 59708 147312 59720 148040
rect 59754 147312 59790 148040
rect 59708 147260 59790 147312
rect 57708 147250 59790 147260
rect 57708 147216 57842 147250
rect 58098 147216 58362 147250
rect 58618 147216 58882 147250
rect 59138 147216 59402 147250
rect 59658 147216 59790 147250
rect 57708 147180 59790 147216
rect 57088 146064 57398 146077
rect 57088 146030 57094 146064
rect 57290 146030 57398 146064
rect 57088 146018 57398 146030
rect 57340 145968 57398 146018
rect 56834 145854 57188 145866
rect 56834 145820 56942 145854
rect 57080 145820 57188 145854
rect 56834 145808 57188 145820
rect 56834 145758 56892 145808
rect 56834 145620 56846 145758
rect 56880 145620 56892 145758
rect 57130 145758 57188 145808
rect 56834 145512 56892 145620
rect 56966 145722 57056 145734
rect 56966 145656 56978 145722
rect 57044 145656 57056 145722
rect 56623 145360 56682 145410
rect 56966 145360 57056 145656
rect 57130 145620 57142 145758
rect 57176 145620 57188 145758
rect 57130 145512 57188 145620
rect 57340 145410 57352 145968
rect 57386 145410 57398 145968
rect 57340 145360 57398 145410
rect 56623 145348 57398 145360
rect 56623 145314 56732 145348
rect 57290 145314 57398 145348
rect 56623 145302 57398 145314
rect 56623 145219 56682 145302
rect 57340 145219 57398 145302
rect 57938 145219 58012 147180
rect 58458 145219 58532 147180
rect 58978 145219 59052 147180
rect 59498 145219 59572 147180
rect 60372 146165 60681 146166
rect 60371 146153 60681 146165
rect 60371 146119 60480 146153
rect 60675 146119 60681 146153
rect 60371 146107 60681 146119
rect 60371 146057 60430 146107
rect 60371 145499 60384 146057
rect 60418 145499 60430 146057
rect 60728 145955 60792 148222
rect 60836 146153 61146 146166
rect 61372 146165 61681 146166
rect 60836 146119 60842 146153
rect 61038 146119 61146 146153
rect 60836 146107 61146 146119
rect 61088 146057 61146 146107
rect 60582 145943 60936 145955
rect 60582 145909 60690 145943
rect 60828 145909 60936 145943
rect 60582 145897 60936 145909
rect 60582 145847 60640 145897
rect 60582 145709 60594 145847
rect 60628 145709 60640 145847
rect 60878 145847 60936 145897
rect 60582 145601 60640 145709
rect 60714 145811 60804 145823
rect 60714 145745 60726 145811
rect 60792 145745 60804 145811
rect 60371 145449 60430 145499
rect 60714 145449 60804 145745
rect 60878 145709 60890 145847
rect 60924 145709 60936 145847
rect 60878 145601 60936 145709
rect 61088 145499 61100 146057
rect 61134 145499 61146 146057
rect 61088 145449 61146 145499
rect 60371 145437 61146 145449
rect 60371 145403 60480 145437
rect 61038 145403 61146 145437
rect 60371 145391 61146 145403
rect 60371 145219 60430 145391
rect 61088 145219 61146 145391
rect 61371 146153 61681 146165
rect 61371 146119 61480 146153
rect 61675 146119 61681 146153
rect 61371 146107 61681 146119
rect 61371 146057 61430 146107
rect 61371 145499 61384 146057
rect 61418 145499 61430 146057
rect 61728 145955 61792 148418
rect 61836 146153 62146 146166
rect 62372 146165 62681 146166
rect 61836 146119 61842 146153
rect 62038 146119 62146 146153
rect 61836 146107 62146 146119
rect 62088 146057 62146 146107
rect 61582 145943 61936 145955
rect 61582 145909 61690 145943
rect 61828 145909 61936 145943
rect 61582 145897 61936 145909
rect 61582 145847 61640 145897
rect 61582 145709 61594 145847
rect 61628 145709 61640 145847
rect 61878 145847 61936 145897
rect 61582 145601 61640 145709
rect 61714 145811 61804 145823
rect 61714 145745 61726 145811
rect 61792 145745 61804 145811
rect 61371 145449 61430 145499
rect 61714 145449 61804 145745
rect 61878 145709 61890 145847
rect 61924 145709 61936 145847
rect 61878 145601 61936 145709
rect 62088 145499 62100 146057
rect 62134 145499 62146 146057
rect 62088 145449 62146 145499
rect 61371 145437 62146 145449
rect 61371 145403 61480 145437
rect 62038 145403 62146 145437
rect 61371 145391 62146 145403
rect 61371 145219 61430 145391
rect 62088 145219 62146 145391
rect 62371 146153 62681 146165
rect 62371 146119 62480 146153
rect 62675 146119 62681 146153
rect 62371 146107 62681 146119
rect 62371 146057 62430 146107
rect 62371 145499 62384 146057
rect 62418 145499 62430 146057
rect 62728 145955 62792 148552
rect 62836 146153 63146 146166
rect 63372 146165 63681 146166
rect 62836 146119 62842 146153
rect 63038 146119 63146 146153
rect 62836 146107 63146 146119
rect 63088 146057 63146 146107
rect 62582 145943 62936 145955
rect 62582 145909 62690 145943
rect 62828 145909 62936 145943
rect 62582 145897 62936 145909
rect 62582 145847 62640 145897
rect 62582 145709 62594 145847
rect 62628 145709 62640 145847
rect 62878 145847 62936 145897
rect 62582 145601 62640 145709
rect 62714 145811 62804 145823
rect 62714 145745 62726 145811
rect 62792 145745 62804 145811
rect 62371 145449 62430 145499
rect 62714 145449 62804 145745
rect 62878 145709 62890 145847
rect 62924 145709 62936 145847
rect 62878 145601 62936 145709
rect 63088 145499 63100 146057
rect 63134 145499 63146 146057
rect 63088 145449 63146 145499
rect 62371 145437 63146 145449
rect 62371 145403 62480 145437
rect 63038 145403 63146 145437
rect 62371 145391 63146 145403
rect 62371 145219 62430 145391
rect 63088 145219 63146 145391
rect 63371 146153 63681 146165
rect 63371 146119 63480 146153
rect 63675 146119 63681 146153
rect 63371 146107 63681 146119
rect 63371 146057 63430 146107
rect 63371 145499 63384 146057
rect 63418 145499 63430 146057
rect 63728 145955 63792 148682
rect 551683 147738 551689 147850
rect 551801 147738 551807 147850
rect 551689 147285 551801 147738
rect 552705 147650 552829 147656
rect 552705 147289 552829 147526
rect 551371 147135 551680 147136
rect 551370 147123 551680 147135
rect 551370 147089 551479 147123
rect 551674 147089 551680 147123
rect 551370 147077 551680 147089
rect 551370 147027 551429 147077
rect 551370 146469 551383 147027
rect 551417 146469 551429 147027
rect 551727 146925 551791 147285
rect 551835 147123 552145 147136
rect 552371 147135 552680 147136
rect 551835 147089 551841 147123
rect 552037 147089 552145 147123
rect 551835 147077 552145 147089
rect 552087 147027 552145 147077
rect 551581 146913 551935 146925
rect 551581 146879 551689 146913
rect 551827 146879 551935 146913
rect 551581 146867 551935 146879
rect 551581 146817 551639 146867
rect 551581 146679 551593 146817
rect 551627 146679 551639 146817
rect 551877 146817 551935 146867
rect 551581 146571 551639 146679
rect 551713 146781 551803 146793
rect 551713 146715 551725 146781
rect 551791 146715 551803 146781
rect 551370 146419 551429 146469
rect 551713 146419 551803 146715
rect 551877 146679 551889 146817
rect 551923 146679 551935 146817
rect 551877 146571 551935 146679
rect 552087 146469 552099 147027
rect 552133 146469 552145 147027
rect 552087 146419 552145 146469
rect 551370 146407 552145 146419
rect 551370 146373 551479 146407
rect 552037 146374 552145 146407
rect 552370 147123 552680 147135
rect 552370 147089 552479 147123
rect 552674 147089 552680 147123
rect 552370 147077 552680 147089
rect 552370 147027 552429 147077
rect 552370 146469 552383 147027
rect 552417 146469 552429 147027
rect 552727 146925 552791 147289
rect 552835 147123 553145 147136
rect 552835 147089 552841 147123
rect 553037 147089 553145 147123
rect 552835 147077 553145 147089
rect 553087 147027 553145 147077
rect 552581 146913 552935 146925
rect 552581 146879 552689 146913
rect 552827 146879 552935 146913
rect 552581 146867 552935 146879
rect 552581 146817 552639 146867
rect 552581 146679 552593 146817
rect 552627 146679 552639 146817
rect 552877 146817 552935 146867
rect 552581 146571 552639 146679
rect 552713 146781 552803 146793
rect 552713 146715 552725 146781
rect 552791 146715 552803 146781
rect 552370 146419 552429 146469
rect 552713 146419 552803 146715
rect 552877 146679 552889 146817
rect 552923 146679 552935 146817
rect 552877 146571 552935 146679
rect 553087 146469 553099 147027
rect 553133 146469 553145 147027
rect 553087 146419 553145 146469
rect 552370 146407 553145 146419
rect 552370 146374 552479 146407
rect 552037 146373 552479 146374
rect 553037 146373 553145 146407
rect 551370 146264 553145 146373
rect 63836 146153 64146 146166
rect 63836 146119 63842 146153
rect 64038 146119 64146 146153
rect 63836 146107 64146 146119
rect 64088 146057 64146 146107
rect 551850 146062 552680 146264
rect 63582 145943 63936 145955
rect 63582 145909 63690 145943
rect 63828 145909 63936 145943
rect 63582 145897 63936 145909
rect 63582 145847 63640 145897
rect 63582 145709 63594 145847
rect 63628 145709 63640 145847
rect 63878 145847 63936 145897
rect 63582 145601 63640 145709
rect 63714 145811 63804 145823
rect 63714 145745 63726 145811
rect 63792 145745 63804 145811
rect 63371 145449 63430 145499
rect 63714 145449 63804 145745
rect 63878 145709 63890 145847
rect 63924 145709 63936 145847
rect 63878 145601 63936 145709
rect 64088 145499 64100 146057
rect 64134 145499 64146 146057
rect 552083 146050 552447 146062
rect 552083 145738 552111 146050
rect 552423 145738 552447 146050
rect 552083 145706 552447 145738
rect 64088 145449 64146 145499
rect 63371 145437 64146 145449
rect 63371 145403 63480 145437
rect 64038 145403 64146 145437
rect 63371 145391 64146 145403
rect 63371 145219 63430 145391
rect 64088 145219 64146 145391
rect 53606 145047 68465 145219
rect 57591 143285 68465 145047
rect 70399 143285 70405 145219
rect 62860 130306 63542 143285
rect 53270 130270 63542 130306
rect 53270 130236 53402 130270
rect 63342 130236 63542 130270
rect 53270 130220 63542 130236
rect 53270 130174 53354 130220
rect 53270 126476 53306 130174
rect 53340 126476 53354 130174
rect 62860 130174 63542 130220
rect 53408 130140 53902 130170
rect 53408 128994 53436 130140
rect 53868 128994 53902 130140
rect 53408 128970 53902 128994
rect 53270 126430 53354 126476
rect 62860 127656 63404 130174
rect 62860 126510 62876 127656
rect 63308 126510 63404 127656
rect 62860 126476 63404 126510
rect 63438 126476 63542 130174
rect 62860 126430 63542 126476
rect 53270 126414 63542 126430
rect 53270 126380 53402 126414
rect 63342 126380 63542 126414
rect 53270 126308 63542 126380
rect 53270 126274 53402 126308
rect 63342 126274 63542 126308
rect 53270 126258 63542 126274
rect 53270 126212 53354 126258
rect 53270 122514 53306 126212
rect 53340 122514 53354 126212
rect 62860 126212 63542 126258
rect 53408 126178 53902 126208
rect 53408 125032 53436 126178
rect 53868 125032 53902 126178
rect 53408 125008 53902 125032
rect 53270 122468 53354 122514
rect 62860 123694 63404 126212
rect 62860 122548 62876 123694
rect 63308 122548 63404 123694
rect 62860 122514 63404 122548
rect 63438 122514 63542 126212
rect 62860 122468 63542 122514
rect 53270 122452 63542 122468
rect 53270 122418 53402 122452
rect 63342 122418 63542 122452
rect 53270 122346 63542 122418
rect 53270 122312 53402 122346
rect 63342 122312 63542 122346
rect 53270 122296 63542 122312
rect 53270 122250 53354 122296
rect 53270 118552 53306 122250
rect 53340 118552 53354 122250
rect 62860 122250 63542 122296
rect 53408 122216 53902 122246
rect 53408 121070 53436 122216
rect 53868 121070 53902 122216
rect 53408 121046 53902 121070
rect 53270 118506 53354 118552
rect 62860 119732 63404 122250
rect 62860 118586 62876 119732
rect 63308 118586 63404 119732
rect 62860 118552 63404 118586
rect 63438 118552 63542 122250
rect 62860 118506 63542 118552
rect 53270 118490 63542 118506
rect 53270 118456 53402 118490
rect 63342 118456 63542 118490
rect 53270 118384 63542 118456
rect 53270 118350 53402 118384
rect 63342 118350 63542 118384
rect 53270 118334 63542 118350
rect 53270 118288 53354 118334
rect 53270 114590 53306 118288
rect 53340 114590 53354 118288
rect 62860 118288 63542 118334
rect 53408 118254 53902 118284
rect 53408 117108 53436 118254
rect 53868 117108 53902 118254
rect 53408 117084 53902 117108
rect 53270 114544 53354 114590
rect 62860 115770 63404 118288
rect 62860 114624 62876 115770
rect 63308 114624 63404 115770
rect 62860 114590 63404 114624
rect 63438 114590 63542 118288
rect 62860 114544 63542 114590
rect 53270 114528 63542 114544
rect 53270 114494 53402 114528
rect 63342 114494 63542 114528
rect 53270 114458 63542 114494
<< rmetal1 >>
rect 60774 150279 61274 150412
<< via1 >>
rect 404827 697923 406599 699695
rect 146520 674731 164088 681965
rect 529691 696526 530082 696917
rect 540137 687119 540399 687288
rect 443952 669616 462134 679662
rect 444062 599950 461834 613648
rect 579580 583476 579810 583706
rect 146784 556095 164076 567969
rect 146694 498073 163458 511617
rect 468092 460100 468156 460164
rect 469092 458614 469156 458678
rect 467592 449422 469659 449507
rect 146500 401839 164068 409147
rect 335668 390738 335732 390802
rect 334668 390082 334732 390146
rect 333824 387884 336416 388772
rect 550243 155065 550317 155139
rect 553806 154223 553982 154275
rect 553713 153977 553765 154195
rect 553816 153897 553992 153949
rect 553817 153581 553993 153633
rect 553713 153335 553765 153553
rect 553815 153255 553991 153307
rect 554354 153333 554406 154316
rect 554659 153337 554711 153581
rect 554967 153333 555019 154316
rect 555269 153334 555325 153578
rect 554410 153236 555264 153288
rect 556092 154372 556536 154425
rect 555954 153331 556006 154318
rect 556050 153331 556102 154318
rect 556146 153331 556198 154318
rect 556242 153331 556294 154318
rect 556338 153331 556390 154318
rect 556434 153331 556486 154318
rect 556530 153331 556582 154318
rect 556019 153226 556436 153278
rect 553786 152694 553867 152746
rect 553690 152448 553742 152666
rect 553787 152367 553868 152419
rect 553788 152053 553869 152105
rect 553690 151806 553742 152024
rect 553787 151725 553868 151777
rect 554277 152768 555439 152820
rect 554226 151746 554278 152722
rect 554520 152349 554583 152728
rect 554834 151741 554886 152717
rect 555135 152348 555198 152727
rect 555446 151741 555498 152717
rect 556266 152772 556416 152824
rect 556197 151742 556249 152727
rect 556293 151740 556345 152727
rect 556397 151742 556449 152727
rect 556223 151644 556294 151696
rect 59229 150309 59303 150383
rect 59506 148852 59570 148916
rect 58986 148640 59050 148704
rect 59644 148682 59708 148746
rect 59114 148552 59178 148616
rect 58462 148464 58526 148528
rect 58590 148418 58654 148482
rect 57942 148292 58006 148356
rect 58078 148222 58142 148286
rect 57928 147988 58010 148042
rect 58058 147392 58110 147968
rect 58448 147988 58530 148042
rect 58578 147392 58630 147968
rect 58968 147988 59050 148042
rect 59098 147392 59150 147968
rect 59488 147988 59570 148042
rect 59618 147392 59670 147968
rect 551689 147738 551801 147850
rect 552705 147526 552829 147650
rect 552111 145738 552423 146050
rect 68465 143285 70399 145219
rect 53436 128994 53868 130140
rect 53436 125032 53868 126178
rect 53436 121070 53868 122216
rect 53436 117108 53868 118254
<< metal2 >>
rect 404827 699695 406599 699701
rect 404818 697923 404827 699695
rect 406599 697923 406608 699695
rect 404827 697917 406599 697923
rect 529662 696917 530093 696928
rect 529662 696526 529691 696917
rect 530082 696526 530093 696917
rect 529662 696509 530093 696526
rect 326218 693564 337501 693970
rect 326218 692489 326803 693564
rect 327878 693559 337501 693564
rect 327878 692494 335984 693559
rect 337049 692494 337501 693559
rect 327878 692489 337501 692494
rect 326218 691947 337501 692489
rect 434817 687328 525966 688544
rect 145394 681965 165394 682901
rect 145394 674731 146520 681965
rect 164088 674731 165394 681965
rect 416733 680130 417949 680139
rect 416733 676381 417949 678914
rect 434817 676381 436033 687328
rect 524750 682605 525966 687328
rect 540110 687288 540426 687322
rect 540110 687119 540137 687288
rect 540399 687119 540426 687288
rect 540110 687092 540426 687119
rect 524750 681389 577407 682605
rect 416733 675165 436033 676381
rect 442918 679662 462918 680730
rect 145394 567969 165394 674731
rect 442918 669616 443952 679662
rect 462134 669616 462918 679662
rect 576191 675517 577407 681389
rect 576187 674311 576196 675517
rect 577402 674311 577411 675517
rect 576191 674306 577407 674311
rect 442918 613648 462918 669616
rect 442918 599950 444062 613648
rect 461834 599950 462918 613648
rect 442918 598730 462918 599950
rect 579559 583706 579826 583727
rect 579559 583476 579580 583706
rect 579810 583476 579826 583706
rect 579559 583451 579826 583476
rect 578155 579543 578375 579547
rect 578150 579538 578380 579543
rect 578150 579318 578155 579538
rect 578375 579318 578380 579538
rect 578150 576166 578380 579318
rect 578150 575927 578380 575936
rect 145394 556095 146784 567969
rect 164076 556095 165394 567969
rect 145394 553901 165394 556095
rect 145398 511617 165398 512901
rect 145398 498073 146694 511617
rect 163458 498073 165398 511617
rect 145398 409147 165398 498073
rect 468083 460100 468092 460164
rect 468156 460100 468165 460164
rect 469083 458614 469092 458678
rect 469156 458614 469165 458678
rect 467580 449507 469674 449521
rect 467580 449422 467592 449507
rect 469659 449422 469674 449507
rect 467580 449411 469674 449422
rect 145398 401839 146500 409147
rect 164068 401839 165398 409147
rect 315391 430218 315511 430227
rect 315391 404023 315407 430218
rect 315496 404023 315511 430218
rect 315391 404007 315511 404023
rect 145398 400903 165398 401839
rect 335657 390802 335741 390811
rect 335657 390738 335668 390802
rect 335732 390738 335741 390802
rect 335657 390728 335741 390738
rect 334650 390146 334758 390164
rect 334650 390082 334668 390146
rect 334732 390082 334758 390146
rect 334650 390066 334758 390082
rect 333727 388772 336528 388853
rect 333727 387884 333824 388772
rect 336416 387884 336528 388772
rect 333727 387811 336528 387884
rect 576858 247713 576970 247718
rect 576854 247611 576863 247713
rect 576965 247611 576974 247713
rect 579976 247705 580088 247710
rect 577650 247697 577762 247702
rect 576858 232630 576970 247611
rect 577646 247595 577655 247697
rect 577757 247595 577766 247697
rect 578446 247661 578558 247666
rect 579244 247661 579356 247666
rect 58562 232518 576970 232630
rect 58044 156733 58160 156746
rect 58044 156631 58049 156733
rect 58151 156631 58160 156733
rect 58044 156620 58160 156631
rect 57942 148356 58006 148365
rect 57933 148292 57942 148348
rect 58006 148292 58015 148348
rect 58052 148292 58126 156620
rect 58462 148528 58526 148537
rect 58462 148455 58526 148464
rect 58572 148488 58646 232518
rect 577650 231478 577762 247595
rect 578442 247559 578451 247661
rect 578553 247559 578562 247661
rect 579240 247559 579249 247661
rect 579351 247559 579360 247661
rect 579972 247603 579981 247705
rect 580083 247603 580092 247705
rect 59080 231366 577762 231478
rect 59092 150383 59166 231366
rect 578446 230244 578558 247559
rect 59584 230132 578558 230244
rect 59612 152171 59686 230132
rect 579244 227180 579356 247559
rect 557468 227068 579356 227180
rect 557468 157815 557580 227068
rect 579976 225946 580088 247603
rect 552845 157703 557580 157815
rect 558758 225834 580088 225946
rect 550237 155065 550243 155139
rect 550317 155065 550323 155139
rect 550243 152171 550317 155065
rect 59612 152097 550317 152171
rect 552845 153073 552957 157703
rect 558758 155853 558870 225834
rect 558758 155732 558870 155741
rect 553794 155321 568284 155379
rect 553794 155207 554446 155321
rect 554560 155207 568284 155321
rect 553794 155179 568284 155207
rect 568484 155179 568493 155379
rect 553794 154275 553994 155179
rect 556256 155073 556320 155179
rect 556256 155000 556320 155009
rect 556086 154425 556542 154431
rect 556086 154422 556092 154425
rect 555614 154372 556092 154422
rect 556536 154372 556542 154425
rect 555614 154366 556542 154372
rect 553794 154223 553806 154275
rect 553982 154223 553994 154275
rect 553794 154217 553994 154223
rect 554348 154316 554411 154327
rect 553707 154195 553771 154201
rect 553707 153977 553713 154195
rect 553765 153977 553771 154195
rect 553707 153553 553771 153977
rect 553804 153949 554004 153956
rect 553804 153897 553816 153949
rect 553992 153897 554004 153949
rect 553804 153891 554004 153897
rect 553861 153831 553994 153891
rect 554348 153831 554354 154316
rect 553861 153698 554354 153831
rect 553861 153640 553994 153698
rect 553804 153633 554004 153640
rect 553804 153581 553817 153633
rect 553993 153581 554004 153633
rect 553804 153575 554004 153581
rect 553707 153335 553713 153553
rect 553765 153335 553771 153553
rect 553707 153073 553771 153335
rect 554348 153333 554354 153698
rect 554406 153831 554411 154316
rect 554961 154316 555024 154327
rect 554961 153831 554967 154316
rect 554406 153698 554967 153831
rect 554406 153333 554411 153698
rect 554348 153327 554411 153333
rect 554650 153581 554721 153590
rect 554650 153337 554659 153581
rect 554715 153337 554721 153581
rect 554650 153327 554721 153337
rect 554961 153333 554967 153698
rect 555019 153333 555024 154316
rect 554961 153327 555024 153333
rect 555259 153578 555335 153590
rect 555259 153334 555269 153578
rect 555325 153334 555335 153578
rect 555259 153325 555335 153334
rect 553803 153307 554003 153313
rect 553803 153255 553815 153307
rect 553991 153255 554003 153307
rect 553803 153248 554003 153255
rect 552845 152961 553771 153073
rect 59229 150383 59303 150389
rect 59092 150309 59229 150383
rect 58986 148704 59050 148713
rect 58986 148631 59050 148640
rect 59092 148616 59166 150309
rect 59229 150303 59303 150309
rect 59506 148916 59570 148925
rect 59506 148843 59570 148852
rect 59612 148752 59686 152097
rect 59612 148746 59708 148752
rect 59612 148682 59644 148746
rect 59612 148676 59708 148682
rect 59092 148552 59114 148616
rect 59178 148552 59184 148616
rect 58572 148482 58654 148488
rect 58572 148418 58590 148482
rect 58572 148412 58654 148418
rect 57942 148283 58006 148292
rect 58052 148286 58142 148292
rect 58052 148222 58078 148286
rect 58052 148216 58142 148222
rect 57916 148044 58024 148054
rect 57916 147988 57928 148044
rect 58010 147988 58024 148044
rect 57916 147978 58024 147988
rect 58052 147968 58126 148216
rect 58436 148044 58544 148054
rect 58436 147988 58448 148044
rect 58530 147988 58544 148044
rect 58436 147978 58544 147988
rect 58052 147392 58058 147968
rect 58110 147392 58126 147968
rect 58052 147376 58126 147392
rect 58572 147968 58646 148412
rect 58956 148044 59064 148054
rect 58956 147988 58968 148044
rect 59050 147988 59064 148044
rect 58956 147978 59064 147988
rect 58572 147392 58578 147968
rect 58630 147392 58646 147968
rect 58572 147376 58646 147392
rect 59092 147968 59166 148552
rect 59476 148044 59584 148054
rect 59476 147988 59488 148044
rect 59570 147988 59584 148044
rect 59476 147978 59584 147988
rect 59092 147392 59098 147968
rect 59150 147392 59166 147968
rect 59092 147376 59166 147392
rect 59612 147968 59686 148676
rect 552845 148177 552957 152961
rect 553684 152957 553771 152961
rect 553870 153099 554003 153248
rect 554404 153288 555272 153294
rect 554404 153236 554410 153288
rect 555264 153236 555272 153288
rect 554404 153230 555272 153236
rect 554764 153099 554897 153230
rect 555614 153099 555747 154366
rect 555948 154318 556010 154325
rect 555948 153761 555954 154318
rect 556006 153761 556010 154318
rect 555948 153406 555951 153761
rect 556007 153406 556010 153761
rect 555948 153331 555954 153406
rect 556006 153331 556010 153406
rect 555948 153325 556010 153331
rect 556044 154318 556106 154325
rect 556044 154261 556050 154318
rect 556102 154261 556106 154318
rect 556044 153906 556047 154261
rect 556103 153906 556106 154261
rect 556044 153331 556050 153906
rect 556102 153331 556106 153906
rect 556044 153325 556106 153331
rect 556140 154318 556202 154325
rect 556140 153761 556146 154318
rect 556198 153761 556202 154318
rect 556140 153406 556143 153761
rect 556199 153406 556202 153761
rect 556140 153331 556146 153406
rect 556198 153331 556202 153406
rect 556140 153325 556202 153331
rect 556236 154318 556298 154325
rect 556236 154261 556242 154318
rect 556294 154261 556298 154318
rect 556236 153906 556239 154261
rect 556295 153906 556298 154261
rect 556236 153331 556242 153906
rect 556294 153331 556298 153906
rect 556236 153325 556298 153331
rect 556332 154318 556394 154325
rect 556332 153761 556338 154318
rect 556390 153761 556394 154318
rect 556332 153406 556335 153761
rect 556391 153406 556394 153761
rect 556332 153331 556338 153406
rect 556390 153331 556394 153406
rect 556332 153325 556394 153331
rect 556428 154318 556490 154325
rect 556428 154261 556434 154318
rect 556486 154261 556490 154318
rect 556428 153906 556431 154261
rect 556487 153906 556490 154261
rect 556428 153331 556434 153906
rect 556486 153331 556490 153906
rect 556428 153325 556490 153331
rect 556524 154318 556586 154325
rect 556524 153761 556530 154318
rect 556582 153853 556586 154318
rect 556623 153906 556679 154261
rect 556582 153761 556915 153853
rect 556524 153406 556527 153761
rect 556583 153729 556915 153761
rect 556583 153406 556586 153729
rect 556524 153331 556530 153406
rect 556582 153331 556586 153406
rect 556524 153325 556586 153331
rect 555996 153278 556446 153284
rect 555996 153226 556019 153278
rect 556436 153226 556446 153278
rect 555996 153220 556446 153226
rect 556163 153099 556296 153220
rect 556791 153155 556915 153729
rect 556791 153141 558879 153155
rect 553870 152966 556415 153099
rect 553684 152666 553748 152957
rect 553870 152904 553951 152966
rect 553797 152826 553951 152904
rect 554748 152826 554881 152966
rect 556282 152855 556415 152966
rect 556163 152845 556415 152855
rect 553797 152756 553875 152826
rect 554272 152820 555446 152826
rect 554272 152768 554277 152820
rect 555439 152768 555446 152820
rect 554272 152762 555446 152768
rect 556163 152778 556178 152845
rect 556271 152830 556415 152845
rect 556791 153039 558763 153141
rect 558865 153039 558879 153141
rect 556791 153031 558879 153039
rect 556271 152824 556432 152830
rect 556163 152772 556266 152778
rect 556416 152772 556432 152824
rect 556163 152766 556432 152772
rect 553779 152746 553875 152756
rect 553779 152694 553786 152746
rect 553867 152694 553875 152746
rect 553779 152688 553875 152694
rect 554214 152722 554282 152734
rect 553684 152448 553690 152666
rect 553742 152448 553748 152666
rect 553684 152024 553748 152448
rect 553779 152419 553876 152426
rect 553779 152367 553787 152419
rect 553868 152367 553876 152419
rect 553779 152358 553876 152367
rect 553799 152258 553876 152358
rect 554214 152258 554226 152722
rect 553799 152181 554226 152258
rect 553799 152114 553876 152181
rect 553780 152105 553876 152114
rect 553780 152053 553788 152105
rect 553869 152053 553876 152105
rect 553780 152046 553876 152053
rect 553684 151806 553690 152024
rect 553742 151806 553748 152024
rect 553684 151799 553748 151806
rect 553780 151777 553876 151785
rect 553780 151725 553787 151777
rect 553868 151725 553876 151777
rect 554214 151746 554226 152181
rect 554278 152258 554282 152722
rect 554502 152728 554593 152734
rect 554502 152725 554520 152728
rect 554502 152341 554516 152725
rect 554583 152349 554593 152728
rect 554581 152341 554593 152349
rect 554502 152329 554593 152341
rect 554824 152717 554892 152734
rect 554824 152258 554834 152717
rect 554278 152181 554834 152258
rect 554278 151746 554282 152181
rect 554214 151734 554282 151746
rect 554824 151741 554834 152181
rect 554886 152258 554892 152717
rect 555119 152727 555216 152734
rect 555119 152724 555135 152727
rect 555198 152724 555216 152727
rect 555119 152335 555130 152724
rect 555206 152335 555216 152724
rect 555119 152325 555216 152335
rect 555438 152717 555506 152734
rect 555438 152258 555446 152717
rect 554886 152181 555446 152258
rect 554886 151741 554892 152181
rect 554824 151734 554892 151741
rect 555438 151741 555446 152181
rect 555498 151741 555506 152717
rect 556192 152727 556255 152734
rect 556192 151884 556197 152727
rect 555438 151734 555506 151741
rect 555990 151788 556197 151884
rect 553780 151257 553876 151725
rect 555990 151257 556086 151788
rect 556192 151742 556197 151788
rect 556249 151742 556255 152727
rect 556192 151734 556255 151742
rect 556289 152727 556350 152734
rect 556289 151740 556293 152727
rect 556345 152687 556350 152727
rect 556349 151844 556350 152687
rect 556345 151740 556350 151844
rect 556289 151734 556350 151740
rect 556392 152727 556454 152734
rect 556392 151742 556397 152727
rect 556449 151742 556454 152727
rect 556555 152656 556693 152665
rect 556791 152656 556915 153031
rect 556555 152532 556564 152656
rect 556688 152532 556915 152656
rect 556555 152523 556693 152532
rect 556189 151696 556302 151702
rect 556189 151633 556200 151696
rect 556294 151644 556302 151696
rect 556283 151633 556302 151644
rect 556189 151625 556302 151633
rect 556392 151257 556472 151742
rect 553780 151161 556472 151257
rect 553780 150962 553876 151161
rect 553780 150857 553876 150866
rect 59612 147392 59618 147968
rect 59670 147392 59686 147968
rect 551689 148065 552957 148177
rect 551689 147850 551801 148065
rect 551689 147732 551801 147738
rect 557740 147650 557864 153031
rect 552699 147526 552705 147650
rect 552829 147526 557864 147650
rect 59612 147376 59686 147392
rect 552083 146050 552447 146078
rect 552083 145738 552111 146050
rect 552423 145738 552447 146050
rect 552083 145706 552447 145738
rect 68465 145219 70399 145225
rect 68461 143290 68465 145214
rect 70399 143290 70403 145214
rect 68465 143279 70399 143285
rect 53408 130140 53902 130170
rect 51537 129678 51639 129682
rect 53408 129678 53436 130140
rect 51532 129673 53436 129678
rect 51532 129571 51537 129673
rect 51639 129571 53436 129673
rect 51532 129566 53436 129571
rect 51537 129562 51639 129566
rect 53408 128994 53436 129566
rect 53868 128994 53902 130140
rect 53408 128970 53902 128994
rect 53408 126178 53902 126208
rect 50987 125538 51089 125542
rect 53408 125538 53436 126178
rect 50982 125533 53436 125538
rect 50982 125431 50987 125533
rect 51089 125431 53436 125533
rect 50982 125426 53436 125431
rect 50987 125422 51089 125426
rect 53408 125032 53436 125426
rect 53868 125032 53902 126178
rect 53408 125008 53902 125032
rect 53408 122216 53902 122246
rect 51653 121604 51755 121608
rect 53408 121604 53436 122216
rect 51648 121599 53436 121604
rect 51648 121497 51653 121599
rect 51755 121497 53436 121599
rect 51648 121492 53436 121497
rect 51653 121488 51755 121492
rect 53408 121070 53436 121492
rect 53868 121070 53902 122216
rect 53408 121046 53902 121070
rect 53408 118254 53902 118284
rect 51487 117418 51589 117422
rect 53408 117418 53436 118254
rect 51482 117413 53436 117418
rect 51482 117311 51487 117413
rect 51589 117311 53436 117413
rect 51482 117306 53436 117311
rect 51487 117302 51589 117306
rect 53408 117108 53436 117306
rect 53868 117108 53902 118254
rect 53408 117084 53902 117108
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 550609 700259 558926 701830
rect 404827 697923 406599 699695
rect 529691 696526 530082 696917
rect 326803 692489 327878 693564
rect 335984 692494 337049 693559
rect 551759 687343 558970 687415
rect 146520 674731 164088 681965
rect 416733 678914 417949 680130
rect 550549 687127 558970 687343
rect 550549 686454 551847 687127
rect 443952 669616 462134 679662
rect 576196 674311 577402 675517
rect 444062 599950 461834 613648
rect 579580 583476 579810 583706
rect 578155 579318 578375 579538
rect 578150 575936 578380 576166
rect 146784 556095 164076 567969
rect 146694 498073 163458 511617
rect 468092 460100 468156 460164
rect 469092 458614 469156 458678
rect 467592 449422 469659 449507
rect 146500 401839 164068 409147
rect 315407 404023 315496 430218
rect 335668 390738 335732 390802
rect 334668 390082 334732 390146
rect 333824 387884 336416 388772
rect 576863 247611 576965 247713
rect 577655 247595 577757 247697
rect 58049 156631 58151 156733
rect 57942 148292 58006 148356
rect 58462 148464 58526 148528
rect 578451 247559 578553 247661
rect 579249 247559 579351 247661
rect 579981 247603 580083 247705
rect 558758 155741 558870 155853
rect 554446 155207 554560 155321
rect 568284 155179 568484 155379
rect 556256 155009 556320 155073
rect 554659 153337 554711 153581
rect 554711 153337 554715 153581
rect 555269 153334 555325 153578
rect 58986 148640 59050 148704
rect 59506 148852 59570 148916
rect 57928 148042 58010 148044
rect 57928 147988 58010 148042
rect 58448 148042 58530 148044
rect 58448 147988 58530 148042
rect 58968 148042 59050 148044
rect 58968 147988 59050 148042
rect 59488 148042 59570 148044
rect 59488 147988 59570 148042
rect 555951 153406 555954 153761
rect 555954 153406 556006 153761
rect 556006 153406 556007 153761
rect 556047 153906 556050 154261
rect 556050 153906 556102 154261
rect 556102 153906 556103 154261
rect 556143 153406 556146 153761
rect 556146 153406 556198 153761
rect 556198 153406 556199 153761
rect 556239 153906 556242 154261
rect 556242 153906 556294 154261
rect 556294 153906 556295 154261
rect 556335 153406 556338 153761
rect 556338 153406 556390 153761
rect 556390 153406 556391 153761
rect 556431 153906 556434 154261
rect 556434 153906 556486 154261
rect 556486 153906 556487 154261
rect 556527 153406 556530 153761
rect 556530 153406 556582 153761
rect 556582 153406 556583 153761
rect 556178 152824 556271 152845
rect 558763 153039 558865 153141
rect 556178 152778 556266 152824
rect 556266 152778 556271 152824
rect 554516 152349 554520 152725
rect 554520 152349 554581 152725
rect 554516 152341 554581 152349
rect 555130 152348 555135 152724
rect 555135 152348 555198 152724
rect 555198 152348 555206 152724
rect 555130 152335 555206 152348
rect 556293 151844 556345 152687
rect 556345 151844 556349 152687
rect 556564 152532 556688 152656
rect 556200 151644 556223 151696
rect 556223 151644 556283 151696
rect 556200 151633 556283 151644
rect 553780 150866 553876 150962
rect 552111 145738 552423 146050
rect 68470 143290 70394 145214
rect 51537 129571 51639 129673
rect 50987 125431 51089 125533
rect 51653 121497 51755 121599
rect 51487 117311 51589 117413
<< metal3 >>
rect 16194 701131 21194 704800
rect 68194 700751 73194 704800
rect 16194 685390 21194 697900
rect 120194 700306 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 68194 693228 73194 697520
rect 120194 695306 196134 700306
rect 68194 688228 182550 693228
rect -800 680242 10218 685242
rect 16194 682901 163994 685390
rect 177550 682901 182550 688228
rect 191134 692480 196134 695306
rect 326798 693564 327883 693569
rect 319829 692489 319835 693564
rect 320910 692489 326803 693564
rect 327878 692489 327883 693564
rect 326798 692484 327883 692489
rect 191134 687480 212060 692480
rect 207060 683876 212060 687480
rect 16194 681965 165394 682901
rect 16194 680390 146520 681965
rect 37396 680389 146520 680390
rect 5218 678990 10218 680242
rect -800 643842 1660 648642
rect -800 633842 1660 638642
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 2546 511946 3024 511957
rect 227 511945 3024 511946
rect 227 511642 2559 511945
rect -800 511530 2559 511642
rect 227 511491 2559 511530
rect 3013 511491 3024 511945
rect 227 511490 3024 511491
rect 2546 511472 3024 511490
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 2022 468600 2504 468610
rect 349 468599 2504 468600
rect 349 468420 2034 468599
rect -800 468308 2034 468420
rect 349 468136 2034 468308
rect 2497 468136 2504 468599
rect 349 468135 2504 468136
rect 2022 468125 2504 468135
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect -800 425086 1694 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 1582 384602 1694 425086
rect 5218 403732 10218 675759
rect 145394 674731 146520 680389
rect 164088 674731 165394 681965
rect 145394 672901 165394 674731
rect 177396 681741 193396 682901
rect 177396 673993 178294 681741
rect 192634 673993 193396 681741
rect 207060 678876 310182 683876
rect 207060 678875 301396 678876
rect 177396 671901 193396 673993
rect 177396 655901 301396 671901
rect 37396 638901 284396 654901
rect 37396 427901 53396 638901
rect 54396 621901 267396 637901
rect 54396 444901 70396 621901
rect 71396 604901 250396 620901
rect 71396 461901 87396 604901
rect 88396 587901 233396 603901
rect 88396 478901 104396 587901
rect 105396 570901 216396 586901
rect 105396 495901 121396 570901
rect 145394 567969 165394 569901
rect 145394 556095 146784 567969
rect 164076 556095 165394 567969
rect 145394 553901 165394 556095
rect 200396 512901 216396 570901
rect 145398 511617 216396 512901
rect 145398 498073 146694 511617
rect 163458 498073 216396 511617
rect 145398 496787 216396 498073
rect 217396 495901 233396 587901
rect 105396 479901 233396 495901
rect 234396 478901 250396 604901
rect 88396 462901 250396 478901
rect 251396 461901 267396 621901
rect 71396 445901 267396 461901
rect 268396 444901 284396 638901
rect 54396 428901 284396 444901
rect 285396 427901 301396 655901
rect 305182 614574 310182 678876
rect 329491 669335 333977 702300
rect 404822 699695 406604 699700
rect 415342 699695 417114 702300
rect 404822 697923 404827 699695
rect 406599 697926 417114 699695
rect 406599 697923 408680 697926
rect 404822 697918 406604 697923
rect 465394 695162 470394 704800
rect 510594 703836 515394 704800
rect 520594 703836 525394 704800
rect 509588 701908 525836 703836
rect 566594 703732 571594 704800
rect 335979 693559 409017 693564
rect 335979 692494 335984 693559
rect 337049 692494 409017 693559
rect 335979 692489 409017 692494
rect 407942 678700 409017 692489
rect 465394 692349 507525 695162
rect 509588 694218 510140 701908
rect 525390 694218 525836 701908
rect 550498 701830 571674 703732
rect 550498 700259 550609 701830
rect 558926 700259 571674 701830
rect 550498 700176 571674 700259
rect 529662 696922 530093 696928
rect 529662 696521 529686 696922
rect 530077 696917 530093 696922
rect 530082 696526 530093 696917
rect 530077 696521 530093 696526
rect 529662 696509 530093 696521
rect 509588 693836 525836 694218
rect 465394 690162 526363 692349
rect 523478 686995 526363 690162
rect 550247 687533 552095 687538
rect 550247 687415 559057 687533
rect 550247 687343 551759 687415
rect 550247 686995 550549 687343
rect 558970 687127 559057 687415
rect 523478 686454 550549 686995
rect 551847 686454 559057 687127
rect 523478 685110 559057 686454
rect 416733 680135 417949 680886
rect 416728 680130 417954 680135
rect 416728 678914 416733 680130
rect 417949 678914 417954 680130
rect 416728 678909 417954 678914
rect 442918 679662 462918 680730
rect 407942 678617 422717 678700
rect 407942 677625 430204 678617
rect 442918 669616 443952 679662
rect 462134 669616 462918 679662
rect 472300 680688 584800 682984
rect 472300 676484 472834 680688
rect 491834 677984 584800 680688
rect 491834 676484 492300 677984
rect 472300 675984 492300 676484
rect 442918 668730 462918 669616
rect 576191 675517 577407 675522
rect 576191 674311 576196 675517
rect 577402 674311 577407 675517
rect 442918 664966 567918 665730
rect 442918 650540 443558 664966
rect 462290 650540 567918 664966
rect 442918 649730 567918 650540
rect 365918 632730 550918 648730
rect 305182 613572 334874 614574
rect 365918 483730 381918 632730
rect 382918 615730 533918 631730
rect 382918 500730 398918 615730
rect 399918 613648 462918 614730
rect 399918 599950 444062 613648
rect 461834 599950 462918 613648
rect 399918 598730 462918 599950
rect 399918 517730 415918 598730
rect 517918 517730 533918 615730
rect 399918 501730 533918 517730
rect 534918 500730 550918 632730
rect 382918 484730 550918 500730
rect 551918 483730 567918 649730
rect 576191 578435 577407 674311
rect 582340 639784 584800 644584
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 579559 583706 579826 583727
rect 578150 583476 579580 583706
rect 579810 583674 583634 583706
rect 579810 583562 584800 583674
rect 579810 583476 583634 583562
rect 578150 579538 578380 583476
rect 579559 583451 579826 583476
rect 578150 579318 578155 579538
rect 578375 579318 578380 579538
rect 578150 579313 578380 579318
rect 576191 577219 580734 578435
rect 578145 576166 578385 576171
rect 578145 575936 578150 576166
rect 578380 575936 578385 576166
rect 578145 575931 578385 575936
rect 365918 467730 567918 483730
rect 578150 460259 578380 575931
rect 579518 560478 580734 577219
rect 579160 555362 583662 560478
rect 579160 550562 584800 555362
rect 579160 545362 583662 550562
rect 579160 544405 584800 545362
rect 579160 543365 579636 544405
rect 580676 543365 584800 544405
rect 579160 540562 584800 543365
rect 579160 540489 583662 540562
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 359782 460164 578380 460259
rect 359782 460100 468092 460164
rect 468156 460100 578380 460164
rect 359782 460029 578380 460100
rect 581011 494252 583774 494348
rect 581011 494140 584800 494252
rect 581011 493920 583774 494140
rect 37396 411901 301396 427901
rect 315391 430218 315511 430227
rect 145398 409147 165398 410903
rect 145398 403732 146500 409147
rect 5218 401839 146500 403732
rect 164068 401839 165398 409147
rect 315391 404023 315407 430218
rect 315496 404023 315511 430218
rect 315391 404007 315511 404023
rect 5218 400903 165398 401839
rect 5218 398732 164798 400903
rect 359782 393971 360012 460029
rect 581011 458843 581439 493920
rect 345229 393741 360012 393971
rect 364943 458678 581439 458843
rect 364943 458614 469092 458678
rect 469156 458614 581439 458678
rect 364943 458415 581439 458614
rect 335668 391085 335732 391091
rect 335668 390811 335732 391021
rect 345229 390883 345459 393741
rect 364943 393188 365371 458415
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 576858 449718 584800 449830
rect 467580 449507 469674 449521
rect 467580 449422 467592 449507
rect 469659 449422 469674 449507
rect 467580 449411 469674 449422
rect 359664 392760 365371 393188
rect 335657 390802 335741 390811
rect 335657 390738 335668 390802
rect 335732 390738 335741 390802
rect 335657 390728 335741 390738
rect 334650 390151 334758 390164
rect 334650 390077 334663 390151
rect 334737 390077 334758 390151
rect 334650 390066 334758 390077
rect 333727 388772 336528 388853
rect 333727 387884 333824 388772
rect 336416 387884 336528 388772
rect 333727 387811 336528 387884
rect 1582 384490 6246 384602
rect -800 381864 4048 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 3936 344426 4048 381864
rect 6134 346444 6246 384490
rect 6134 346332 24260 346444
rect 3936 344314 19792 344426
rect -800 338642 15754 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect -800 295420 7532 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 7420 260508 7532 295420
rect 15642 268318 15754 338642
rect 19680 272558 19792 344314
rect 24148 275304 24260 346332
rect 24148 275192 38092 275304
rect 19680 272446 34188 272558
rect 15642 268206 30922 268318
rect 7420 260396 19588 260508
rect -800 252398 13750 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 13638 149840 13750 252398
rect 19476 151614 19588 260396
rect 30810 153354 30922 268206
rect 34076 154942 34188 272446
rect 37980 156738 38092 275192
rect 576858 247713 576970 449718
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 576858 247611 576863 247713
rect 576965 247611 576970 247713
rect 576858 247606 576970 247611
rect 577650 405296 584800 405408
rect 577650 247697 577762 405296
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 577650 247595 577655 247697
rect 577757 247595 577762 247697
rect 577650 247590 577762 247595
rect 578446 358874 584800 358986
rect 578446 247661 578558 358874
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 578446 247559 578451 247661
rect 578553 247559 578558 247661
rect 578446 247554 578558 247559
rect 579244 313652 584800 313764
rect 579244 247661 579356 313652
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 579244 247559 579249 247661
rect 579351 247559 579356 247661
rect 579976 269230 584800 269342
rect 579976 247705 580088 269230
rect 579976 247603 579981 247705
rect 580083 247603 580088 247705
rect 579976 247598 580088 247603
rect 579244 247554 579356 247559
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 582378 202438 583422 225230
rect 570134 201394 583422 202438
rect 37980 156733 58156 156738
rect 37980 156631 58049 156733
rect 58151 156631 58156 156733
rect 37980 156626 58156 156631
rect 558753 155853 558875 155858
rect 558753 155741 558758 155853
rect 558870 155741 558875 155853
rect 558753 155736 558875 155741
rect 554441 155321 554565 155326
rect 554441 155207 554446 155321
rect 554560 155207 554565 155321
rect 34076 154830 59604 154942
rect 30810 153242 59072 153354
rect 19476 151502 58554 151614
rect 13638 149728 58040 149840
rect 57928 148356 58040 149728
rect 57928 148292 57942 148356
rect 58006 148292 58040 148356
rect 57928 148092 58040 148292
rect 57920 148054 58040 148092
rect 58442 148528 58554 151502
rect 58442 148464 58462 148528
rect 58526 148464 58554 148528
rect 58442 148076 58554 148464
rect 58960 148704 59072 153242
rect 58960 148640 58986 148704
rect 59050 148640 59072 148704
rect 58960 148076 59072 148640
rect 59492 148916 59604 154830
rect 554441 152734 554565 155207
rect 556251 155073 556325 155078
rect 556251 155009 556256 155073
rect 556320 155009 556325 155073
rect 556251 155004 556325 155009
rect 556256 154266 556320 155004
rect 556042 154261 556108 154266
rect 556042 153906 556047 154261
rect 556103 154179 556108 154261
rect 556234 154261 556320 154266
rect 556234 154179 556239 154261
rect 556103 153995 556239 154179
rect 556103 153906 556108 153995
rect 556042 153901 556108 153906
rect 556234 153906 556239 153995
rect 556295 154179 556320 154261
rect 556426 154261 556492 154266
rect 556426 154179 556431 154261
rect 556295 153995 556431 154179
rect 556295 153906 556300 153995
rect 556234 153901 556300 153906
rect 556426 153906 556431 153995
rect 556487 153906 556492 154261
rect 556426 153901 556492 153906
rect 555946 153761 556012 153766
rect 554650 153581 554721 153590
rect 554650 153337 554659 153581
rect 554715 153460 554721 153581
rect 555259 153578 555335 153590
rect 555259 153460 555269 153578
rect 554715 153390 555269 153460
rect 554715 153337 554721 153390
rect 554650 153327 554721 153337
rect 555259 153334 555269 153390
rect 555325 153460 555335 153578
rect 555325 153334 555362 153460
rect 555946 153406 555951 153761
rect 556007 153679 556012 153761
rect 556138 153761 556204 153766
rect 556138 153679 556143 153761
rect 556007 153495 556143 153679
rect 556007 153406 556012 153495
rect 555946 153401 556012 153406
rect 556138 153406 556143 153495
rect 556199 153679 556204 153761
rect 556330 153761 556396 153766
rect 556330 153679 556335 153761
rect 556199 153495 556335 153679
rect 556199 153406 556204 153495
rect 556138 153401 556204 153406
rect 556330 153406 556335 153495
rect 556391 153679 556396 153761
rect 556522 153761 556588 153766
rect 556522 153679 556527 153761
rect 556391 153495 556527 153679
rect 556391 153406 556396 153495
rect 556330 153401 556396 153406
rect 556522 153406 556527 153495
rect 556583 153406 556588 153761
rect 556522 153401 556588 153406
rect 555259 153325 555362 153334
rect 554441 152725 554593 152734
rect 554441 152516 554516 152725
rect 554502 152341 554516 152516
rect 554581 152640 554593 152725
rect 555119 152724 555216 152734
rect 555119 152640 555130 152724
rect 554581 152516 555130 152640
rect 554581 152341 554593 152516
rect 554502 152329 554593 152341
rect 555119 152335 555130 152516
rect 555206 152335 555216 152724
rect 555119 152325 555216 152335
rect 553775 150962 553881 150967
rect 553775 150866 553780 150962
rect 553876 150866 553881 150962
rect 553775 150861 553881 150866
rect 59492 148852 59506 148916
rect 59570 148852 59604 148916
rect 59492 148110 59604 148852
rect 59488 148076 59604 148110
rect 58440 148054 58560 148076
rect 58960 148054 59080 148076
rect 59480 148054 59604 148076
rect 57916 148044 58040 148054
rect 57916 147988 57928 148044
rect 58010 147988 58040 148044
rect 57916 147982 58040 147988
rect 58436 148044 58560 148054
rect 58436 147988 58448 148044
rect 58530 147988 58560 148044
rect 58436 147982 58560 147988
rect 58956 148044 59080 148054
rect 58956 147988 58968 148044
rect 59050 147988 59080 148044
rect 58956 147982 59080 147988
rect 59476 148044 59604 148054
rect 59476 147988 59488 148044
rect 59570 147988 59604 148044
rect 59476 147986 59604 147988
rect 553780 150689 553876 150861
rect 555292 150689 555362 153325
rect 558758 153141 558870 155736
rect 568279 155379 568489 155384
rect 570134 155379 571178 201394
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect 568279 155179 568284 155379
rect 568484 155179 571178 155379
rect 568279 155174 568489 155179
rect 558758 153039 558763 153141
rect 558865 153039 558870 153141
rect 558758 153034 558870 153039
rect 556163 152845 556287 152855
rect 556163 152778 556178 152845
rect 556271 152778 556287 152845
rect 556163 152766 556287 152778
rect 556164 151706 556225 152766
rect 556288 152692 556350 152701
rect 556288 152687 556354 152692
rect 556288 151844 556293 152687
rect 556349 152656 556354 152687
rect 556559 152656 556693 152661
rect 556349 152532 556564 152656
rect 556688 152532 556693 152656
rect 556349 151844 556354 152532
rect 556559 152527 556693 152532
rect 556288 151834 556354 151844
rect 556164 151696 556302 151706
rect 556164 151633 556200 151696
rect 556283 151633 556302 151696
rect 556164 151616 556302 151633
rect 553780 150593 555362 150689
rect 59476 147982 59600 147986
rect 57916 147978 58024 147982
rect 58436 147978 58544 147982
rect 58956 147978 59064 147982
rect 59476 147978 59584 147982
rect 552106 146050 552428 146055
rect 552106 145738 552111 146050
rect 552423 145738 552428 146050
rect 552106 145733 552428 145738
rect 552111 145219 552423 145733
rect 553780 145219 553876 150593
rect 582340 146830 584800 151630
rect 68465 145214 583122 145219
rect 68465 143290 68470 145214
rect 70394 143290 583122 145214
rect 68465 143285 583122 143290
rect 581188 141630 583122 143285
rect 581188 138734 584800 141630
rect 582340 136830 584800 138734
rect 30464 129673 51644 129678
rect 30464 129571 51537 129673
rect 51639 129571 51644 129673
rect 30464 129566 51644 129571
rect 30464 124888 30576 129566
rect -800 124776 30576 124888
rect 34286 125533 51094 125538
rect 34286 125431 50987 125533
rect 51089 125431 51094 125533
rect 34286 125426 51094 125431
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 34286 81666 34398 125426
rect -800 81554 34398 81666
rect 39560 121599 51760 121604
rect 39560 121497 51653 121599
rect 51755 121497 51760 121599
rect 39560 121492 51760 121497
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 39560 38444 39672 121492
rect -800 38332 39672 38444
rect 46468 117413 51594 117418
rect 46468 117311 51487 117413
rect 51589 117311 51594 117413
rect 46468 117306 51594 117311
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 46468 17022 46580 117306
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 46580 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< rmetal3 >>
rect 15291 697900 21689 701131
rect 67397 697520 73795 700751
rect 4490 675759 10888 678990
<< via3 >>
rect 319835 692489 320910 693564
rect 2559 511491 3013 511945
rect 2034 468136 2497 468599
rect 146520 674731 164088 681965
rect 178294 673993 192634 681741
rect 146784 556095 164076 567969
rect 510140 694218 525390 701908
rect 529686 696917 530077 696922
rect 529686 696526 529691 696917
rect 529691 696526 530077 696917
rect 529686 696521 530077 696526
rect 443952 669616 462134 679662
rect 472834 676484 491834 680688
rect 329310 625656 329890 666846
rect 443558 650540 462290 664966
rect 327010 615420 327590 625656
rect 579636 543365 580676 544405
rect 146500 401839 164068 409147
rect 315407 404023 315496 430218
rect 335668 391021 335732 391085
rect 467592 449422 469659 449507
rect 334663 390146 334737 390151
rect 334663 390082 334668 390146
rect 334668 390082 334732 390146
rect 334732 390082 334737 390146
rect 334663 390077 334737 390082
rect 333824 387884 336416 388772
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702908 222294 704800
rect 227594 702908 232594 704800
rect 318994 703328 323994 704800
rect 329294 703328 334294 704800
rect 217076 694329 313018 702908
rect 318994 702300 334294 703328
rect 319734 701870 333977 702300
rect 509588 702016 525836 702728
rect 217076 694064 326008 694329
rect 303443 693564 326008 694064
rect 303443 692489 319835 693564
rect 320910 692489 326008 693564
rect 303443 685915 326008 692489
rect 145394 681965 165394 682901
rect 145394 674731 146520 681965
rect 164088 674731 165394 681965
rect 145394 672901 165394 674731
rect 177396 681741 193396 682901
rect 177396 673993 178294 681741
rect 192634 673993 193396 681741
rect 177396 672901 193396 673993
rect 37396 655903 301396 671903
rect 318008 668449 326008 685915
rect 329491 680766 333977 701870
rect 344882 701908 525836 702016
rect 344882 694218 510140 701908
rect 525390 696917 525836 701908
rect 529662 696922 530093 696928
rect 529662 696917 529686 696922
rect 525390 696526 529686 696917
rect 525390 694218 525836 696526
rect 529662 696521 529686 696526
rect 530077 696521 530093 696922
rect 529662 696509 530093 696521
rect 344882 694016 525836 694218
rect 329491 669335 333996 680766
rect 344882 679466 352882 694016
rect 509588 693836 525836 694016
rect 419347 680730 454676 683321
rect 419347 680128 462918 680730
rect 344618 671466 352882 679466
rect 318008 667405 326803 668449
rect 318008 666882 329224 667405
rect 318008 666856 329488 666882
rect 318008 666846 329900 666856
rect 2546 511945 3024 511957
rect 2546 511491 2559 511945
rect 3013 511491 3024 511945
rect 2546 511472 3024 511491
rect 2022 468599 2504 468610
rect 2022 468136 2034 468599
rect 2497 468136 2504 468599
rect 2022 468125 2504 468136
rect 37396 427903 53396 655903
rect 54394 638901 284394 654901
rect 54394 444901 70394 638901
rect 71394 621901 267394 637901
rect 71394 461901 87394 621901
rect 88394 604901 250394 620901
rect 88394 478901 104394 604901
rect 105394 587901 233394 604017
rect 105394 495901 121394 587901
rect 122394 567969 165394 569901
rect 122394 556095 146784 567969
rect 164076 556095 165394 567969
rect 122394 553901 165394 556095
rect 122394 512901 138394 553901
rect 217394 512901 233394 587901
rect 122394 496901 233394 512901
rect 234394 495901 250394 604901
rect 105394 479901 250394 495901
rect 251394 478901 267394 621901
rect 88394 462901 267394 478901
rect 268394 461901 284394 638901
rect 71394 445901 284394 461901
rect 285394 444901 301394 655903
rect 318008 641449 329310 666846
rect 320810 625656 329310 641449
rect 329890 625656 329900 666846
rect 333349 625826 333996 669335
rect 344882 650788 352882 671466
rect 442918 679662 462918 680128
rect 442918 669616 443952 679662
rect 462134 669616 462918 679662
rect 472300 680688 492300 680984
rect 472300 676484 472834 680688
rect 491834 676484 492300 680688
rect 472300 675984 492300 676484
rect 442918 668730 462918 669616
rect 365918 664966 462918 665730
rect 365918 650540 443558 664966
rect 462290 650540 462918 664966
rect 365918 649730 462918 650540
rect 320810 625646 327010 625656
rect 327000 615420 327010 625646
rect 327590 625646 329900 625656
rect 327590 615420 327600 625646
rect 327000 615410 327600 615420
rect 355680 594766 356922 618535
rect 345203 593524 356922 594766
rect 345203 453097 346445 593524
rect 365918 483730 381918 649730
rect 382918 632730 567918 648730
rect 382918 500730 398918 632730
rect 399918 615730 550918 631730
rect 399918 517730 415918 615730
rect 470918 613524 533918 614730
rect 470918 599798 472272 613524
rect 489906 599798 533918 613524
rect 470918 598730 533918 599798
rect 517918 517730 533918 598730
rect 399918 501730 533918 517730
rect 534918 500730 550918 615730
rect 382918 484730 550918 500730
rect 551918 483730 567918 632730
rect 579635 544405 580677 544406
rect 579635 543365 579636 544405
rect 580676 543365 580677 544405
rect 579635 543364 580677 543365
rect 365918 467730 567918 483730
rect 350636 460921 385103 460945
rect 350636 455969 350660 460921
rect 355612 456299 385103 460921
rect 355612 455969 380103 456299
rect 350636 455945 380103 455969
rect 345203 451855 364263 453097
rect 363221 449507 364263 451855
rect 467580 449507 469674 449521
rect 363221 449422 467592 449507
rect 469659 449422 484266 449507
rect 363221 448557 484266 449422
rect 363841 445744 484266 448557
rect 54394 428901 301394 444901
rect 315391 430218 315711 430227
rect 37396 411903 165398 427903
rect 145398 409147 165398 411903
rect 145398 401839 146500 409147
rect 164068 401839 165398 409147
rect 315391 404023 315407 430218
rect 315644 404023 315711 430218
rect 315391 404007 315711 404023
rect 145398 400903 165398 401839
rect 363221 388853 364263 390887
rect 333727 388772 364263 388853
rect 333727 387884 333824 388772
rect 336416 387884 364263 388772
rect 333727 387811 364263 387884
<< via4 >>
rect 146520 674731 164088 681965
rect 178294 673993 192634 681741
rect 510140 694218 525390 701908
rect 2582 511514 2990 511922
rect 2057 468159 2474 468576
rect 146784 556095 164076 567969
rect 329310 625656 329890 666846
rect 443952 669616 462134 679662
rect 472834 676484 491834 680688
rect 327010 615420 327590 625656
rect 472272 599798 489906 613524
rect 579659 543388 580653 544382
rect 350660 455969 355612 460921
rect 380103 451299 385103 456299
rect 146500 401839 164068 409147
rect 315407 404023 315496 430218
rect 315496 404023 315644 430218
rect 335540 391085 335860 391213
rect 335540 391021 335668 391085
rect 335668 391021 335732 391085
rect 335732 391021 335860 391085
rect 335540 390893 335860 391021
rect 334540 390151 334860 390274
rect 334540 390077 334663 390151
rect 334663 390077 334737 390151
rect 334737 390077 334860 390151
rect 334540 389954 334860 390077
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 703568 180894 704800
rect 175894 702568 200140 703568
rect 217294 702908 222294 704800
rect 227594 702908 232594 704800
rect 318994 703328 323994 704800
rect 329294 703328 334294 704800
rect 175894 702300 180894 702568
rect 199140 694994 200140 702568
rect 199140 693994 215608 694994
rect 217076 694329 313018 702908
rect 318994 702300 334294 703328
rect 319734 701870 333977 702300
rect 509588 702016 525836 702728
rect 217076 694064 326008 694329
rect 214608 686056 215608 693994
rect 303443 685915 326008 694064
rect 145394 681965 165394 682901
rect 145394 674731 146520 681965
rect 164088 674731 165394 681965
rect 145394 672901 165394 674731
rect 177396 681741 193396 682901
rect 177396 673993 178294 681741
rect 192634 673993 193396 681741
rect 177396 672901 193396 673993
rect 37396 655903 301396 671903
rect 318008 668449 326008 685915
rect 329491 680766 333977 701870
rect 344882 701908 525836 702016
rect 344882 694218 510140 701908
rect 525390 694218 525836 701908
rect 344882 694016 525836 694218
rect 329491 669335 333996 680766
rect 344882 679466 352882 694016
rect 422585 692424 428028 694016
rect 509588 693836 525836 694016
rect 419347 680730 454676 683321
rect 472300 680730 492300 680984
rect 419347 680128 462918 680730
rect 344618 671466 352882 679466
rect 318008 667405 326803 668449
rect 318008 667076 329224 667405
rect 318008 666846 330218 667076
rect 2546 511946 3024 511957
rect 2546 511922 8768 511946
rect 2546 511514 2582 511922
rect 2990 511514 8768 511922
rect 2546 511490 8768 511514
rect 2546 511472 3024 511490
rect 2022 468600 2504 468610
rect 2022 468576 7099 468600
rect 2022 468159 2057 468576
rect 2474 468159 7099 468576
rect 2022 468135 7099 468159
rect 2022 468125 2504 468135
rect 6634 390402 7099 468135
rect 8312 391482 8768 511490
rect 37396 427903 53396 655903
rect 54394 638901 284394 654901
rect 54394 444901 70394 638901
rect 71394 621901 267394 637901
rect 71394 461901 87394 621901
rect 88394 604901 250394 620901
rect 88394 478901 104394 604901
rect 105394 587901 233394 604017
rect 105394 495901 121394 587901
rect 122394 567969 165394 569901
rect 122394 556095 146784 567969
rect 164076 556095 165394 567969
rect 122394 553901 165394 556095
rect 122394 512901 138394 553901
rect 217394 512901 233394 587901
rect 122394 496901 233394 512901
rect 234394 495901 250394 604901
rect 105394 479901 250394 495901
rect 251394 478901 267394 621901
rect 88394 462901 267394 478901
rect 268394 461901 284394 638901
rect 71394 445901 284394 461901
rect 285394 444901 301394 655903
rect 318008 641449 329310 666846
rect 320810 625656 329310 641449
rect 329890 625656 330218 666846
rect 333349 625826 333996 669335
rect 344882 650788 352882 671466
rect 442918 679662 462918 680128
rect 442918 669616 443952 679662
rect 462134 669616 462918 679662
rect 442918 668730 462918 669616
rect 470918 680688 492300 680730
rect 470918 676484 472834 680688
rect 491834 676484 492300 680688
rect 470918 675984 492300 676484
rect 470918 665730 490918 675984
rect 470918 649730 567918 665730
rect 365918 632730 550918 648730
rect 320810 615420 327010 625656
rect 327590 625550 330218 625656
rect 327590 615420 327934 625550
rect 320810 614586 327934 615420
rect 320810 595474 325810 614586
rect 320810 590474 338214 595474
rect 333214 460945 338214 590474
rect 365918 483730 381918 632730
rect 382918 615730 533918 631730
rect 382918 500730 398918 615730
rect 399918 613524 490918 614730
rect 399918 599798 472272 613524
rect 489906 599798 490918 613524
rect 399918 598730 490918 599798
rect 399918 517730 415918 598730
rect 517918 517730 533918 615730
rect 399918 501730 533918 517730
rect 534918 500730 550918 632730
rect 382918 484730 550918 500730
rect 551918 483730 567918 649730
rect 365918 467730 567918 483730
rect 579635 544382 580677 544406
rect 579635 543388 579659 544382
rect 580653 543388 580677 544382
rect 333214 460921 355636 460945
rect 333214 455969 350660 460921
rect 355612 455969 355636 460921
rect 579635 459210 580677 543388
rect 333214 455945 355636 455969
rect 361201 458168 580677 459210
rect 333214 454104 338214 455945
rect 54394 428901 301394 444901
rect 315381 453776 338214 454104
rect 315381 453774 332876 453776
rect 315381 430218 315711 453774
rect 361201 448109 362243 458168
rect 380079 456299 385127 456323
rect 380079 451299 380103 456299
rect 385103 451299 385127 456299
rect 380079 451275 385127 451299
rect 380103 450246 385103 451275
rect 380103 445246 411181 450246
rect 37396 411903 165398 427903
rect 145398 409147 165398 411903
rect 145398 401839 146500 409147
rect 164068 401839 165398 409147
rect 315381 404023 315407 430218
rect 315644 404023 315711 430218
rect 315381 403997 315711 404023
rect 145398 400903 165398 401839
rect 8312 391213 338981 391482
rect 8312 391026 335540 391213
rect 335516 390893 335540 391026
rect 335860 391026 338981 391213
rect 335860 390893 335884 391026
rect 335516 390869 335884 390893
rect 339620 390402 340085 392808
rect 6634 390274 340085 390402
rect 6634 389954 334540 390274
rect 334860 389954 340085 390274
rect 6634 389937 340085 389954
rect 334516 389930 334884 389937
rect 258138 281192 274538 281592
rect 256138 280792 276938 281192
rect 254538 280392 278538 280792
rect 252138 279992 264538 280392
rect 269338 279992 280938 280392
rect 250138 279592 258938 279992
rect 274138 279592 282538 279992
rect 248938 279192 256538 279592
rect 276538 279192 283738 279592
rect 247338 278792 253738 279192
rect 278938 278792 285338 279192
rect 246538 278392 252538 278792
rect 261338 278392 261738 278792
rect 262538 278392 271338 278792
rect 272138 278392 272538 278792
rect 280538 278392 286538 278792
rect 245738 277992 250938 278392
rect 258938 277992 273338 278392
rect 273738 277992 274538 278392
rect 282138 277992 287338 278392
rect 244538 277592 249338 277992
rect 255738 277592 277338 277992
rect 283738 277592 288538 277992
rect 243338 277192 248538 277592
rect 253738 277192 262138 277592
rect 262538 277192 263738 277592
rect 268538 277192 268938 277592
rect 269738 277192 279738 277592
rect 284938 277192 289738 277592
rect 242538 276792 247338 277192
rect 253338 276792 258538 277192
rect 259338 276792 259738 277192
rect 273338 276792 280538 277192
rect 286138 276792 290538 277192
rect 241338 276392 245738 276792
rect 250538 276392 256538 276792
rect 276938 276392 282138 276792
rect 287338 276392 291338 276792
rect 240538 275992 244938 276392
rect 249738 275992 254538 276392
rect 278538 275992 283738 276392
rect 288138 275992 292138 276392
rect 240138 275592 244138 275992
rect 248538 275592 252938 275992
rect 280538 275592 284138 275992
rect 289338 275592 292938 275992
rect 238938 275192 242938 275592
rect 246938 275192 250938 275592
rect 282138 275192 285738 275592
rect 290538 275192 293738 275592
rect 238138 274792 242138 275192
rect 246138 274792 249738 275192
rect 282938 274792 287338 275192
rect 290938 274792 294538 275192
rect 237738 274392 241338 274792
rect 244938 274392 248938 274792
rect 284138 274392 287738 274792
rect 291738 274392 294938 274792
rect 236938 273992 240138 274392
rect 244538 273992 247738 274392
rect 285738 273992 289338 274392
rect 292938 273992 295738 274392
rect 236138 273592 239738 273992
rect 243338 273592 246138 273992
rect 286538 273592 290138 273992
rect 293738 273592 296538 273992
rect 235738 273192 238938 273592
rect 242938 273192 245738 273592
rect 287738 273192 290538 273592
rect 294138 273192 296938 273592
rect 234938 272792 238138 273192
rect 241338 272792 244538 273192
rect 288938 272792 292138 273192
rect 295338 272792 297738 273192
rect 234138 272392 237338 272792
rect 240538 272392 243738 272792
rect 289338 272392 292538 272792
rect 295738 272392 298538 272792
rect 233738 271992 236938 272392
rect 239738 271992 242938 272392
rect 264938 271992 265738 272392
rect 290538 271992 292938 272392
rect 296538 271992 298938 272392
rect 232938 271592 236138 271992
rect 239338 271592 241338 271992
rect 259738 271592 262138 271992
rect 232538 271192 235338 271592
rect 238538 271192 241338 271592
rect 258538 271192 262138 271592
rect 231738 270792 234938 271192
rect 237738 270792 240538 271192
rect 257338 270792 262138 271192
rect 231338 270392 234138 270792
rect 236938 270392 239738 270792
rect 254938 270392 262138 270792
rect 262938 270792 264138 271992
rect 264938 271592 271738 271992
rect 272538 271592 274138 271992
rect 291338 271592 294138 271992
rect 297338 271592 299738 271992
rect 264538 271192 275338 271592
rect 292138 271192 294538 271592
rect 298138 271192 300538 271592
rect 264538 270792 276538 271192
rect 292538 270792 295338 271192
rect 298538 270792 300938 271192
rect 262938 270392 263738 270792
rect 264938 270392 266138 270792
rect 230538 269992 233338 270392
rect 236538 269992 238938 270392
rect 254138 269992 263338 270392
rect 264138 269992 265338 270392
rect 230138 269592 232938 269992
rect 236138 269592 238138 269992
rect 253338 269592 259338 269992
rect 229738 269192 232138 269592
rect 235338 269192 237738 269592
rect 252138 269192 259338 269592
rect 228938 268792 231738 269192
rect 234538 268792 236938 269192
rect 251738 268792 259338 269192
rect 228538 268392 231338 268792
rect 234138 268392 236538 268792
rect 250538 268392 259338 268792
rect 261738 268792 265338 269992
rect 266938 269592 268538 270792
rect 270138 270392 276938 270792
rect 277338 270392 278538 270792
rect 293738 270392 295738 270792
rect 299338 270392 301338 270792
rect 268938 269992 269738 270392
rect 270938 269992 271338 270392
rect 272138 269992 279738 270392
rect 294138 269992 296938 270392
rect 299738 269992 302138 270392
rect 268938 269592 270138 269992
rect 273738 269592 280538 269992
rect 294938 269592 297338 269992
rect 300138 269592 302538 269992
rect 266938 269192 271338 269592
rect 272138 269192 273338 269592
rect 274138 269192 282538 269592
rect 295338 269192 297738 269592
rect 300938 269192 302938 269592
rect 261738 268392 264938 268792
rect 266938 268392 269738 269192
rect 270138 268392 271338 269192
rect 271738 268792 273738 269192
rect 274138 268792 282938 269192
rect 296138 268792 298538 269192
rect 301338 268792 303738 269192
rect 272138 268392 284138 268792
rect 296938 268392 298938 268792
rect 302138 268392 304138 268792
rect 228138 267992 230538 268392
rect 233338 267992 235338 268392
rect 249738 267992 253338 268392
rect 256138 267992 259338 268392
rect 260938 267992 262138 268392
rect 227738 267592 230138 267992
rect 232938 267592 234938 267992
rect 248938 267592 254538 267992
rect 256538 267592 262138 267992
rect 262938 267592 264138 268392
rect 265338 267992 269338 268392
rect 272138 267992 273338 268392
rect 273738 267992 284538 268392
rect 297338 267992 299738 268392
rect 302538 267992 304538 268392
rect 265338 267592 270938 267992
rect 271338 267592 273338 267992
rect 274538 267592 275738 267992
rect 227338 267192 229738 267592
rect 232538 267192 234538 267592
rect 248138 267192 254938 267592
rect 256538 267192 258138 267592
rect 258538 267192 264538 267592
rect 226938 266792 229338 267192
rect 231738 266792 233738 267192
rect 247338 266792 252138 267192
rect 252538 266792 254938 267192
rect 226538 266392 228938 266792
rect 231338 266392 233338 266792
rect 226138 265992 228538 266392
rect 230538 265992 232938 266392
rect 246138 265992 251738 266792
rect 252938 266392 254938 266792
rect 255738 266792 264538 267192
rect 265338 267192 273338 267592
rect 276138 267192 280938 267992
rect 281338 267592 286138 267992
rect 298138 267592 300138 267992
rect 302938 267592 305338 267992
rect 282938 267192 286538 267592
rect 298538 267192 300538 267592
rect 303338 267192 305738 267592
rect 265338 266792 266938 267192
rect 267338 266792 273338 267192
rect 255738 266392 258538 266792
rect 259738 266392 262138 266792
rect 262938 266392 264538 266792
rect 265738 266392 266138 266792
rect 267338 266392 268538 266792
rect 268938 266392 273338 266792
rect 274138 266392 277338 267192
rect 277738 266792 281338 267192
rect 282138 266792 283338 267192
rect 284138 266792 286938 267192
rect 298938 266792 301338 267192
rect 303738 266792 306138 267192
rect 277738 266392 281738 266792
rect 282138 266392 283738 266792
rect 284538 266392 288138 266792
rect 299738 266392 301738 266792
rect 304538 266392 306538 266792
rect 225338 265592 227738 265992
rect 230538 265592 232138 265992
rect 245338 265592 251738 265992
rect 224938 265192 227338 265592
rect 230138 265192 231738 265592
rect 244938 265192 251738 265592
rect 224538 264792 226938 265192
rect 229338 264792 231338 265192
rect 244538 264792 248138 265192
rect 248538 264792 251738 265192
rect 253338 265992 257338 266392
rect 260538 265992 262138 266392
rect 263738 265992 264938 266392
rect 266538 265992 268138 266392
rect 269338 265992 269738 266392
rect 271738 265992 272938 266392
rect 274138 265992 279338 266392
rect 280138 265992 284138 266392
rect 284938 265992 289338 266392
rect 300138 265992 302138 266392
rect 304938 265992 306938 266392
rect 253338 265592 256938 265992
rect 253338 264792 255338 265592
rect 255738 265192 256938 265592
rect 258938 265192 260138 265592
rect 260938 265192 262538 265992
rect 256138 264792 257338 265192
rect 224138 264392 226538 264792
rect 228938 264392 230538 264792
rect 244138 264392 250538 264792
rect 251338 264392 252538 264792
rect 253738 264392 254938 264792
rect 255738 264392 257338 264792
rect 258538 264792 262538 265192
rect 262938 264792 265338 265992
rect 266538 265592 268538 265992
rect 268938 265592 270138 265992
rect 266138 265192 270138 265592
rect 266138 264792 267738 265192
rect 268538 264792 270138 265192
rect 271738 265592 273338 265992
rect 276138 265592 279338 265992
rect 279738 265592 280938 265992
rect 282138 265592 285738 265992
rect 286538 265592 289738 265992
rect 300938 265592 302938 265992
rect 305338 265592 307338 265992
rect 271738 265192 274138 265592
rect 258538 264392 262138 264792
rect 268938 264392 269738 264792
rect 271738 264392 274538 265192
rect 277338 264792 280938 265592
rect 282538 265192 286138 265592
rect 286938 265192 290538 265592
rect 301338 265192 302938 265592
rect 305738 265192 307738 265592
rect 281738 264792 282138 265192
rect 283738 264792 286538 265192
rect 287338 264792 291338 265192
rect 301738 264792 303338 265192
rect 306138 264792 308138 265192
rect 276138 264392 278538 264792
rect 278938 264392 287738 264792
rect 288138 264392 291738 264792
rect 302138 264392 304138 264792
rect 306538 264392 308538 264792
rect 223738 263992 226138 264392
rect 228538 263992 230538 264392
rect 243738 263992 246938 264392
rect 247338 263992 250938 264392
rect 251338 263992 252938 264392
rect 223338 263592 225738 263992
rect 228138 263592 230138 263992
rect 243338 263592 246538 263992
rect 247338 263592 249338 263992
rect 250138 263592 251738 263992
rect 252138 263592 252938 263992
rect 254138 263592 257738 264392
rect 258538 263992 260538 264392
rect 261338 263992 261738 264392
rect 272538 263992 274138 264392
rect 276138 263992 278138 264392
rect 278938 263992 285338 264392
rect 286138 263992 287738 264392
rect 289338 263992 292138 264392
rect 302938 263992 304538 264392
rect 306938 263992 308938 264392
rect 258938 263592 260138 263992
rect 276138 263592 279738 263992
rect 280538 263592 284538 263992
rect 286538 263592 288138 263992
rect 289338 263592 292538 263992
rect 303338 263592 304938 263992
rect 307338 263592 309338 263992
rect 222938 263192 225338 263592
rect 227738 263192 229338 263592
rect 242938 263192 249738 263592
rect 250138 263192 251338 263592
rect 252538 263192 253338 263592
rect 254138 263192 257338 263592
rect 276138 263192 281338 263592
rect 282538 263192 285738 263592
rect 286938 263192 288138 263592
rect 290138 263192 292538 263592
rect 303738 263192 305738 263592
rect 307738 263192 309738 263592
rect 222538 262792 224938 263192
rect 227338 262792 228938 263192
rect 242538 262792 248138 263192
rect 248538 262792 249738 263192
rect 250538 262792 250938 263192
rect 222138 262392 224538 262792
rect 226538 262392 228538 262792
rect 241338 262392 247738 262792
rect 248538 262392 250138 262792
rect 252138 262392 253738 263192
rect 254138 262792 255738 263192
rect 276938 262792 281738 263192
rect 282938 262792 286138 263192
rect 288538 262792 289738 263192
rect 290538 262792 293738 263192
rect 304138 262792 305738 263192
rect 308138 262792 310138 263192
rect 254538 262392 255338 262792
rect 278138 262392 278938 262792
rect 279738 262392 282538 262792
rect 284138 262392 286138 262792
rect 222138 261992 224138 262392
rect 226538 261992 228138 262392
rect 241338 261992 242938 262392
rect 243338 261992 244538 262392
rect 244938 261992 247338 262392
rect 248938 261992 250138 262392
rect 250938 261992 253738 262392
rect 279738 261992 282938 262392
rect 284538 261992 286138 262392
rect 221738 261592 223738 261992
rect 226138 261592 227738 261992
rect 240938 261592 242538 261992
rect 221338 261192 223338 261592
rect 225738 261192 227338 261592
rect 240538 261192 242538 261592
rect 243338 261592 246538 261992
rect 248938 261592 253338 261992
rect 280138 261592 284138 261992
rect 284938 261592 286138 261992
rect 288138 262392 290138 262792
rect 288138 261992 290538 262392
rect 291738 261992 294138 262792
rect 304538 262392 306138 262792
rect 308538 262392 310538 262792
rect 304938 261992 306938 262392
rect 308938 261992 310938 262392
rect 288138 261592 290138 261992
rect 290938 261592 294538 261992
rect 305338 261592 306938 261992
rect 309338 261592 311338 261992
rect 243338 261192 244938 261592
rect 249338 261192 252138 261592
rect 281738 261192 284538 261592
rect 220938 260792 222938 261192
rect 225338 260792 226938 261192
rect 239738 260792 242138 261192
rect 242938 260792 244938 261192
rect 245738 260792 247338 261192
rect 248938 260792 251738 261192
rect 282538 260792 284538 261192
rect 284938 261192 286538 261592
rect 286938 261192 287738 261592
rect 288938 261192 289338 261592
rect 284938 260792 288138 261192
rect 290538 260792 292538 261592
rect 292938 260792 294938 261592
rect 305738 261192 307338 261592
rect 309738 261192 311738 261592
rect 306138 260792 308138 261192
rect 310138 260792 312138 261192
rect 220538 260392 222538 260792
rect 224938 260392 226538 260792
rect 239338 260392 241738 260792
rect 242538 260392 244538 260792
rect 245338 260392 247738 260792
rect 248138 260392 251338 260792
rect 282938 260392 284538 260792
rect 285338 260392 288138 260792
rect 289738 260392 295738 260792
rect 306538 260392 308538 260792
rect 310538 260392 312538 260792
rect 220138 259992 222138 260392
rect 224538 259992 226138 260392
rect 238938 259992 241738 260392
rect 242138 259992 244138 260392
rect 245338 259992 250138 260392
rect 283338 259992 284138 260392
rect 284938 259992 288138 260392
rect 219738 259592 222138 259992
rect 224138 259592 225738 259992
rect 238538 259592 243738 259992
rect 219738 259192 221738 259592
rect 223738 259192 225338 259592
rect 237738 259192 243738 259592
rect 245738 259592 246938 259992
rect 247338 259592 250138 259992
rect 284538 259592 288138 259992
rect 245738 259192 248938 259592
rect 284538 259192 286938 259592
rect 287338 259192 288138 259592
rect 288938 259992 296138 260392
rect 306938 259992 308538 260392
rect 310938 259992 312938 260392
rect 288938 259592 290538 259992
rect 291338 259592 293738 259992
rect 294138 259592 296938 259992
rect 307338 259592 308938 259992
rect 288938 259192 290938 259592
rect 291338 259192 297338 259592
rect 307738 259192 309338 259592
rect 311338 259192 313338 259992
rect 219338 258792 221338 259192
rect 223738 258792 224938 259192
rect 237338 258792 244138 259192
rect 245738 258792 248538 259192
rect 284938 258792 286938 259192
rect 288538 258792 292138 259192
rect 292938 258792 294538 259192
rect 295338 258792 297338 259192
rect 308138 258792 309738 259192
rect 311738 258792 313738 259192
rect 218938 258392 220938 258792
rect 222938 258392 224538 258792
rect 236938 258392 239738 258792
rect 240138 258392 242138 258792
rect 218538 257992 220538 258392
rect 218538 257592 220138 257992
rect 222538 257592 224138 258392
rect 236938 257992 239338 258392
rect 240138 257992 241738 258392
rect 242538 257992 244538 258792
rect 245338 258392 247738 258792
rect 288138 258392 289338 258792
rect 245338 257992 247338 258392
rect 236538 257592 239738 257992
rect 242938 257592 244138 257992
rect 245738 257592 247338 257992
rect 287738 257992 289338 258392
rect 290138 258392 292138 258792
rect 293338 258392 294938 258792
rect 295738 258392 297738 258792
rect 308538 258392 309738 258792
rect 312138 258392 314138 258792
rect 290138 257992 292538 258392
rect 293338 257992 298138 258392
rect 308938 257992 310538 258392
rect 312538 257992 314538 258392
rect 287738 257592 289738 257992
rect 290138 257592 292938 257992
rect 218138 257192 219738 257592
rect 222138 257192 223738 257592
rect 236138 257192 240138 257592
rect 246138 257192 246538 257592
rect 287738 257192 293338 257592
rect 294138 257192 296138 257992
rect 217738 256792 219738 257192
rect 221738 256792 223338 257192
rect 235738 256792 240138 257192
rect 243338 256792 244138 257192
rect 288538 256792 291338 257192
rect 217338 256392 219338 256792
rect 217338 255992 218938 256392
rect 221338 255992 222938 256792
rect 235738 256392 237738 256792
rect 234938 255992 237338 256392
rect 238138 255992 239738 256792
rect 240538 256392 241738 256792
rect 242938 256392 244538 256792
rect 216938 255592 218938 255992
rect 220938 255592 222538 255992
rect 234938 255592 237738 255992
rect 238538 255592 239338 255992
rect 240138 255592 241738 256392
rect 242538 255592 244538 256392
rect 289338 256392 291338 256792
rect 291738 256792 293338 257192
rect 291738 256392 292938 256792
rect 294538 256392 296138 257192
rect 296538 257192 298538 257992
rect 309338 257192 310938 257992
rect 312938 257592 314938 257992
rect 313338 257192 314938 257592
rect 296538 256792 298938 257192
rect 309738 256792 311338 257192
rect 313338 256792 315338 257192
rect 297338 256392 299338 256792
rect 310138 256392 311738 256792
rect 313738 256392 315738 256792
rect 289338 255992 292538 256392
rect 289738 255592 292538 255992
rect 293338 255592 294938 256392
rect 297338 255992 299738 256392
rect 297738 255592 299738 255992
rect 310538 255592 312138 256392
rect 314138 255992 316138 256392
rect 314538 255592 316138 255992
rect 216538 255192 218538 255592
rect 220538 255192 222138 255592
rect 216538 254792 218138 255192
rect 216138 254392 218138 254792
rect 220138 254392 221738 255192
rect 234538 254792 238138 255592
rect 240138 255192 241338 255592
rect 242538 255192 244138 255592
rect 240538 254792 241738 255192
rect 242938 254792 244138 255192
rect 290538 254792 292138 255592
rect 292938 255192 295338 255592
rect 298138 255192 300138 255592
rect 310938 255192 312538 255592
rect 314538 255192 316538 255592
rect 293338 254792 295738 255192
rect 234538 254392 236138 254792
rect 237338 254392 239738 254792
rect 240538 254392 242138 254792
rect 260938 254392 272938 254792
rect 290938 254392 292938 254792
rect 293738 254392 296138 254792
rect 296938 254392 300538 255192
rect 311338 254792 312938 255192
rect 314938 254792 316938 255192
rect 215738 253992 217738 254392
rect 219738 253992 221338 254392
rect 233738 253992 235738 254392
rect 215738 253592 217338 253992
rect 215338 253192 217338 253592
rect 219338 253592 220938 253992
rect 233338 253592 235738 253992
rect 238138 253992 240138 254392
rect 240538 253992 241738 254392
rect 260538 253992 273738 254392
rect 238138 253592 241738 253992
rect 259738 253592 274938 253992
rect 291738 253592 293338 254392
rect 294138 253992 296138 254392
rect 296538 253992 298538 254392
rect 294138 253592 298138 253992
rect 298938 253592 300938 254392
rect 311738 253992 313338 254792
rect 315338 254392 316938 254792
rect 315338 253992 317338 254392
rect 312138 253592 313738 253992
rect 315738 253592 317338 253992
rect 219338 253192 220538 253592
rect 233338 253192 236138 253592
rect 237338 253192 241738 253592
rect 257338 253192 276138 253592
rect 292138 253192 301338 253592
rect 312538 253192 314138 253592
rect 214938 252792 216938 253192
rect 218938 252792 220538 253192
rect 232938 252792 241738 253192
rect 256538 252792 276538 253192
rect 292538 252792 294538 253192
rect 214938 252392 216538 252792
rect 214538 251992 216538 252392
rect 218538 252392 220138 252792
rect 218538 251992 219738 252392
rect 232538 251992 234138 252792
rect 234538 252392 238938 252792
rect 239738 252392 241738 252792
rect 255738 252392 270138 252792
rect 270938 252392 277738 252792
rect 234538 251992 236538 252392
rect 237338 251992 241338 252392
rect 255738 251992 263738 252392
rect 264538 251992 270138 252392
rect 271338 251992 278138 252392
rect 214538 251592 216138 251992
rect 218138 251592 219738 251992
rect 232138 251592 236538 251992
rect 238538 251592 240538 251992
rect 255338 251592 262938 251992
rect 266138 251592 269738 251992
rect 214138 251192 215738 251592
rect 218138 251192 219338 251592
rect 232138 251192 237738 251592
rect 213738 250792 215738 251192
rect 217738 250792 218938 251192
rect 231738 250792 235338 251192
rect 213738 250392 215338 250792
rect 217338 250392 218938 250792
rect 213338 249592 214938 250392
rect 217338 249992 218538 250392
rect 216938 249592 218138 249992
rect 212938 249192 214938 249592
rect 216538 249192 218138 249592
rect 231338 249192 232938 250792
rect 233338 249992 235338 250792
rect 236138 250392 237738 251192
rect 238938 250792 240538 251592
rect 254938 251192 262938 251592
rect 265338 251192 265738 251592
rect 254538 250792 258138 251192
rect 258538 250792 260538 251192
rect 253338 250392 257738 250792
rect 236138 249992 238938 250392
rect 252538 249992 257338 250392
rect 258538 249992 260138 250792
rect 261338 250392 262938 251192
rect 264938 250392 266138 251192
rect 266938 250792 269738 251592
rect 270938 251592 278538 251992
rect 292938 251592 294538 252792
rect 295338 251992 296938 253192
rect 295738 251592 296938 251992
rect 297738 252792 301338 253192
rect 312938 252792 314138 253192
rect 316138 253192 317738 253592
rect 316138 252792 318138 253192
rect 297738 251992 302138 252792
rect 312938 252392 314538 252792
rect 316538 252392 318138 252792
rect 313338 251992 314938 252392
rect 297738 251592 300138 251992
rect 300538 251592 302138 251992
rect 313738 251592 314938 251992
rect 316938 251992 318538 252392
rect 316938 251592 318938 251992
rect 270938 251192 272538 251592
rect 273338 251192 279338 251592
rect 233738 249592 237338 249992
rect 212938 248792 214538 249192
rect 216538 248792 217738 249192
rect 230938 248792 232938 249192
rect 234538 248792 236938 249592
rect 237738 249192 238938 249992
rect 252138 249592 256938 249992
rect 252138 249192 256538 249592
rect 257738 249192 260138 249992
rect 260938 249992 263338 250392
rect 260938 249592 263738 249992
rect 264938 249592 266538 250392
rect 260938 249192 266538 249592
rect 238138 248792 238538 249192
rect 251738 248792 256538 249192
rect 212538 247992 214138 248792
rect 216138 248392 217738 248792
rect 216138 247992 217338 248392
rect 230538 247992 232538 248792
rect 234938 248392 237338 248792
rect 251338 248392 256538 248792
rect 257338 248792 260138 249192
rect 260538 248792 266538 249192
rect 267338 248792 269338 250792
rect 270538 250392 272538 251192
rect 270138 249992 272538 250392
rect 269738 249592 272538 249992
rect 273738 250792 280138 251192
rect 273738 250392 275738 250792
rect 276938 250392 280538 250792
rect 293738 250392 295338 251592
rect 296138 251192 297338 251592
rect 298138 251192 299738 251592
rect 300538 251192 302938 251592
rect 313738 251192 315338 251592
rect 296138 250392 297738 251192
rect 273738 249992 275338 250392
rect 277338 249992 280938 250392
rect 294538 249992 295738 250392
rect 296538 249992 297738 250392
rect 298938 250792 300138 251192
rect 301338 250792 302938 251192
rect 314138 250792 315338 251192
rect 317338 251192 318938 251592
rect 317338 250792 319338 251192
rect 298938 249992 300538 250792
rect 301338 249992 303338 250792
rect 273738 249592 274938 249992
rect 275738 249592 276538 249992
rect 277738 249592 281338 249992
rect 269738 249192 272138 249592
rect 236138 247992 238138 248392
rect 250938 247992 256138 248392
rect 212138 247192 213738 247992
rect 215738 247192 216938 247992
rect 230538 247592 233738 247992
rect 234538 247592 238138 247992
rect 250538 247592 256138 247992
rect 211738 246392 213338 247192
rect 215338 246792 216938 247192
rect 230138 247192 238138 247592
rect 250138 247192 253338 247592
rect 230138 246792 237738 247192
rect 249738 246792 252938 247192
rect 253738 246792 256138 247592
rect 215338 246392 216538 246792
rect 229738 246392 237338 246792
rect 211338 245592 212938 246392
rect 210938 244792 212538 245592
rect 214938 245192 216138 246392
rect 229738 245592 231338 246392
rect 232138 245992 237338 246392
rect 249338 245992 252538 246792
rect 253338 245992 256138 246792
rect 257338 247992 269738 248792
rect 257338 247192 262538 247992
rect 263338 247592 270138 247992
rect 270938 247592 272138 249192
rect 263338 247192 268538 247592
rect 268938 247192 270538 247592
rect 271338 247192 272138 247592
rect 273338 249192 274938 249592
rect 273338 247192 274538 249192
rect 275338 248792 276938 249592
rect 278138 249192 281738 249592
rect 294938 249192 296138 249992
rect 296938 249592 297738 249992
rect 299338 249592 303338 249992
rect 314538 250392 315738 250792
rect 317738 250392 319338 250792
rect 314538 249592 316138 250392
rect 318138 249592 319738 250392
rect 275338 247992 276538 248792
rect 278538 248392 282538 249192
rect 295338 248792 297338 249192
rect 298538 248792 298938 249192
rect 299738 248792 303738 249592
rect 314938 249192 316538 249592
rect 318138 249192 320138 249592
rect 278138 247992 282938 248392
rect 295738 247992 304138 248792
rect 315338 248392 316938 249192
rect 318538 248792 320538 249192
rect 275338 247192 276938 247992
rect 278138 247592 279338 247992
rect 277738 247192 279338 247592
rect 280138 247192 283338 247992
rect 257338 246792 262138 247192
rect 263338 246792 268138 247192
rect 269338 246792 270938 247192
rect 273338 246792 274938 247192
rect 257338 245992 261338 246792
rect 262938 246392 268138 246792
rect 269738 246392 270938 246792
rect 273738 246392 274938 246792
rect 275338 246392 279738 247192
rect 262938 245992 265338 246392
rect 228938 245192 232538 245592
rect 214538 244792 215738 245192
rect 210538 244392 212538 244792
rect 210538 243592 212138 244392
rect 214138 243992 215738 244792
rect 228938 244792 232938 245192
rect 233338 244792 237338 245992
rect 248938 245592 252138 245992
rect 252938 245592 256538 245992
rect 248938 245192 256538 245592
rect 257738 245192 261338 245992
rect 262538 245592 265338 245992
rect 265738 245992 268538 246392
rect 269738 245992 270538 246392
rect 265738 245592 269338 245992
rect 273338 245592 279738 246392
rect 262138 245192 265338 245592
rect 266138 245192 270138 245592
rect 248538 244792 256938 245192
rect 257738 244792 259338 245192
rect 228938 244392 236938 244792
rect 248138 244392 259338 244792
rect 218138 243992 219338 244392
rect 228938 243992 230538 244392
rect 230938 243992 234938 244392
rect 247338 243992 252138 244392
rect 253738 243992 258938 244392
rect 210138 243192 212138 243592
rect 213738 243192 215338 243992
rect 217738 243592 219338 243992
rect 210138 242392 211738 243192
rect 213738 242792 214938 243192
rect 209738 241192 211338 242392
rect 213338 241992 214938 242792
rect 217338 242792 218938 243592
rect 228538 243192 230538 243992
rect 231338 243592 234538 243992
rect 231738 243192 234538 243592
rect 246938 243592 252138 243992
rect 254138 243592 258938 243992
rect 259738 243992 261338 245192
rect 261738 244792 265738 245192
rect 261738 244392 263338 244792
rect 264138 244392 265738 244792
rect 266538 244792 270538 245192
rect 272938 244792 279738 245592
rect 266538 244392 271738 244792
rect 246938 243192 251738 243592
rect 254538 243192 258538 243592
rect 220138 242792 221338 243192
rect 217338 242392 221338 242792
rect 228138 242792 230538 243192
rect 234938 242792 236138 243192
rect 228138 242392 233338 242792
rect 217738 241992 220938 242392
rect 213338 241592 214538 241992
rect 218138 241592 220538 241992
rect 228138 241592 233738 242392
rect 234538 241992 236138 242792
rect 246538 242792 251738 243192
rect 252138 242792 254138 243192
rect 234938 241592 235738 241992
rect 246538 241592 254138 242792
rect 254938 241992 256138 243192
rect 212938 241192 214138 241592
rect 209338 240392 210938 241192
rect 208938 239592 210938 240392
rect 212538 239992 214138 241192
rect 228138 240792 230138 241592
rect 230538 241192 233738 241592
rect 246538 241192 250938 241592
rect 231338 240792 231738 241192
rect 232138 240792 233338 241192
rect 228138 240392 229738 240792
rect 232138 240392 232538 240792
rect 246538 240392 248938 241192
rect 249738 240392 250938 241192
rect 251338 241192 254138 241592
rect 254538 241192 256538 241992
rect 251338 240392 256938 241192
rect 257338 240792 258538 243192
rect 259738 242792 260938 243992
rect 261738 243592 262938 244392
rect 264138 243592 266138 244392
rect 261738 243192 263338 243592
rect 262138 242792 263738 243192
rect 264538 242792 266138 243592
rect 266938 243592 271338 244392
rect 272938 243992 274138 244792
rect 272538 243592 274138 243992
rect 266938 243192 268538 243592
rect 267338 242792 268538 243192
rect 259338 242392 261338 242792
rect 262138 242392 264138 242792
rect 259338 241992 261738 242392
rect 262538 241992 264138 242392
rect 264538 241992 266538 242792
rect 259338 241592 264138 241992
rect 264938 241592 266538 241992
rect 267338 242392 268938 242792
rect 269338 242392 271338 243592
rect 272138 243192 274138 243592
rect 271738 242792 274138 243192
rect 274938 243592 279738 244792
rect 280538 246792 283738 247192
rect 296138 246792 300138 247992
rect 300538 247592 304538 247992
rect 315738 247592 316938 248392
rect 318938 247992 320538 248792
rect 300938 247192 304538 247592
rect 300538 246792 304538 247192
rect 316138 247192 317338 247592
rect 319338 247192 320938 247992
rect 316138 246792 317738 247192
rect 280538 246392 284138 246792
rect 296138 246392 297738 246792
rect 299338 246392 300138 246792
rect 300938 246392 302538 246792
rect 280538 245992 284538 246392
rect 296138 245992 297338 246392
rect 299338 245992 300538 246392
rect 280538 245592 284938 245992
rect 280538 244392 282138 245592
rect 282538 244792 285338 245592
rect 297338 245192 298138 245592
rect 298938 245192 300538 245992
rect 296938 244792 298538 245192
rect 299338 244792 300538 245192
rect 301338 245992 302538 246392
rect 302938 245992 304938 246792
rect 316538 246392 317738 246792
rect 319738 246392 321338 247192
rect 316538 245992 318138 246392
rect 301338 245592 304938 245992
rect 316938 245592 318138 245992
rect 320138 245592 321738 246392
rect 301338 244792 305338 245592
rect 316938 245192 318538 245592
rect 280138 243992 282138 244392
rect 280138 243592 281738 243992
rect 282938 243592 285738 244792
rect 296938 244392 298938 244792
rect 300138 244392 305338 244792
rect 317338 244792 318538 245192
rect 320538 245192 321738 245592
rect 317338 244392 318938 244792
rect 320538 244392 322138 245192
rect 296938 243992 298538 244392
rect 300138 243992 302138 244392
rect 303738 243992 305338 244392
rect 317738 243992 318938 244392
rect 297338 243592 299338 243992
rect 300138 243592 301738 243992
rect 302538 243592 305738 243992
rect 317738 243592 319338 243992
rect 320938 243592 322538 244392
rect 271738 242392 273738 242792
rect 274938 242392 278138 243592
rect 267338 241592 271338 242392
rect 259338 241192 264538 241592
rect 259738 240792 264538 241192
rect 265338 241192 266538 241592
rect 267738 241192 271738 241592
rect 272138 241192 273738 242392
rect 274538 241992 278138 242392
rect 278538 241992 281738 243592
rect 282538 243192 285738 243592
rect 298138 243192 301338 243592
rect 302138 243192 305738 243592
rect 282538 242792 286138 243192
rect 298138 242792 300138 243192
rect 282538 242392 286538 242792
rect 274538 241592 281738 241992
rect 257338 240392 259338 240792
rect 259738 240392 261338 240792
rect 261738 240392 264938 240792
rect 228138 239992 230138 240392
rect 230538 239992 230938 240392
rect 231738 239992 234538 240392
rect 212538 239592 213738 239992
rect 219338 239592 220538 239992
rect 208938 238792 210538 239592
rect 212138 238792 213738 239592
rect 218938 239192 220938 239592
rect 208538 237592 210138 238792
rect 212138 237992 213338 238792
rect 218538 238392 221338 239192
rect 228138 238792 234938 239992
rect 218138 237992 221738 238392
rect 227738 237992 229338 238792
rect 229738 238392 234938 238792
rect 229738 237992 232938 238392
rect 233338 237992 234938 238392
rect 246538 239192 248538 240392
rect 249738 239592 256938 240392
rect 257738 239992 260938 240392
rect 262138 239992 264938 240392
rect 265338 239992 266938 241192
rect 269338 240792 273738 241192
rect 274938 240792 281738 241592
rect 282138 241192 286538 242392
rect 298538 241992 300138 242792
rect 300938 242392 306138 243192
rect 318138 242792 319338 243592
rect 321338 242792 322938 243592
rect 298938 241592 300138 241992
rect 300538 241992 306138 242392
rect 318538 241992 319738 242792
rect 321738 241992 322938 242792
rect 300538 241592 302538 241992
rect 304138 241592 306538 241992
rect 298938 241192 302538 241592
rect 270138 240392 274138 240792
rect 267738 239992 268538 240392
rect 270138 239992 274538 240392
rect 274938 239992 281338 240792
rect 282138 239992 286938 241192
rect 298538 240792 302538 241192
rect 304538 240792 306538 241592
rect 318538 241192 320138 241992
rect 321738 241592 323338 241992
rect 318938 240792 320138 241192
rect 322138 241192 323338 241592
rect 298938 239992 302538 240792
rect 303338 239992 304138 240392
rect 304938 239992 306538 240792
rect 257738 239592 260538 239992
rect 262538 239592 266938 239992
rect 267338 239592 268938 239992
rect 249338 239192 257338 239592
rect 257738 239192 260938 239592
rect 262938 239192 268938 239592
rect 269738 239192 280538 239992
rect 282138 239592 286538 239992
rect 298938 239592 300938 239992
rect 281738 239192 286538 239592
rect 246538 238792 261738 239192
rect 262938 238792 279338 239192
rect 246538 238392 279338 238792
rect 279738 238792 280938 239192
rect 281338 238792 286538 239192
rect 246538 237992 255338 238392
rect 256138 237992 278938 238392
rect 208138 236792 210138 237592
rect 208138 235992 209738 236792
rect 211738 236392 212938 237992
rect 218138 237192 219738 237992
rect 217738 236392 219338 237192
rect 211738 235992 212538 236392
rect 207738 235192 209738 235992
rect 207738 233992 209338 235192
rect 211338 234792 212538 235992
rect 217738 235592 219738 236392
rect 220138 235592 221738 237992
rect 227338 237192 229338 237992
rect 230938 237592 232938 237992
rect 231338 237192 232938 237592
rect 246538 237192 254938 237992
rect 256538 237592 278938 237992
rect 279738 237992 283338 238792
rect 284138 237992 286538 238792
rect 256938 237192 262938 237592
rect 227738 236792 230538 237192
rect 231338 236792 234538 237192
rect 246538 236792 248538 237192
rect 248938 236792 254538 237192
rect 257738 236792 259338 237192
rect 260538 236792 262938 237192
rect 227738 236392 234538 236792
rect 227338 235992 234938 236392
rect 211338 234392 212138 234792
rect 217738 234392 221738 235592
rect 210938 233992 212138 234392
rect 207338 233592 209338 233992
rect 207338 232392 208938 233592
rect 210538 233192 212138 233992
rect 218138 233992 221738 234392
rect 226938 235592 232538 235992
rect 232938 235592 234938 235992
rect 246138 235992 248538 236792
rect 249338 236392 254138 236792
rect 258138 236392 259338 236792
rect 261338 236392 262938 236792
rect 248938 235992 253738 236392
rect 261738 235992 262938 236392
rect 264138 236792 266138 237592
rect 267338 237192 272538 237592
rect 273338 237192 279338 237592
rect 279738 237192 282938 237992
rect 283738 237592 286538 237992
rect 299338 239192 300138 239592
rect 299338 238792 300538 239192
rect 299338 238392 300938 238792
rect 301338 238392 302538 239992
rect 302938 239592 304538 239992
rect 304938 239592 306938 239992
rect 312538 239592 314138 239992
rect 302938 238792 306938 239592
rect 312138 238792 314538 239592
rect 319338 239192 320538 240792
rect 322138 240392 323738 241192
rect 322538 239192 324138 240392
rect 319738 238792 320938 239192
rect 299338 237992 302538 238392
rect 299338 237592 300938 237992
rect 267338 236792 269338 237192
rect 271738 236792 272538 237192
rect 274138 236792 282938 237192
rect 283338 236792 286538 237592
rect 299738 237192 300938 237592
rect 301338 237592 302538 237992
rect 303338 237592 306938 238792
rect 301338 237192 304938 237592
rect 305338 237192 306538 237592
rect 264138 236392 265738 236792
rect 267738 236392 268938 236792
rect 274138 236392 286138 236792
rect 264138 235992 265338 236392
rect 267738 235992 268138 236392
rect 274538 235992 286138 236392
rect 218138 233592 221338 233992
rect 218538 233192 221338 233592
rect 210938 232792 211738 233192
rect 218538 232792 220938 233192
rect 206938 230792 208938 232392
rect 210538 231592 211738 232792
rect 218938 232392 220938 232792
rect 226938 232392 228938 235592
rect 229738 235192 230538 235592
rect 230938 235192 232538 235592
rect 233338 235192 234538 235592
rect 230938 234792 232938 235192
rect 229738 234392 232938 234792
rect 229338 233992 232938 234392
rect 229338 233592 232538 233992
rect 229338 233192 232938 233592
rect 233338 233192 234538 233592
rect 229738 232792 230538 233192
rect 230938 232392 234938 233192
rect 246138 232792 248138 235992
rect 248938 235592 252538 235992
rect 264538 235592 264938 235992
rect 275338 235592 276938 235992
rect 277338 235592 278538 235992
rect 279338 235592 286138 235992
rect 248938 235192 251738 235592
rect 275738 235192 276138 235592
rect 277738 235192 278538 235592
rect 248938 234792 251338 235192
rect 279738 234792 286138 235592
rect 299738 235192 300538 237192
rect 301338 236792 306538 237192
rect 312538 236792 314538 238792
rect 315738 237592 316938 238792
rect 319738 237992 321338 238792
rect 315338 237192 316938 237592
rect 320138 237192 321338 237992
rect 322938 238392 324138 239192
rect 322938 237592 324538 238392
rect 323338 237192 324538 237592
rect 315338 236792 317338 237192
rect 320138 236792 321738 237192
rect 301338 235192 302538 236792
rect 302938 236392 306538 236792
rect 311738 236392 317338 236792
rect 303338 235592 306938 236392
rect 311338 235992 317338 236392
rect 310938 235592 317338 235992
rect 302938 235192 306938 235592
rect 248938 233192 250938 234792
rect 280138 234392 286538 234792
rect 280138 233992 282938 234392
rect 280538 233592 282938 233992
rect 283338 233592 286538 234392
rect 299338 234392 300938 235192
rect 301338 234792 306938 235192
rect 299338 233992 300538 234392
rect 301738 233992 302538 234792
rect 302938 234392 306938 234792
rect 310538 235192 317338 235592
rect 310538 234392 312138 235192
rect 312538 234792 314538 235192
rect 315338 234792 317338 235192
rect 303338 233992 306938 234392
rect 248538 232792 250538 233192
rect 219738 231992 220138 232392
rect 226538 231992 228938 232392
rect 229338 231992 230138 232392
rect 214938 231592 216138 231992
rect 226538 231592 230538 231992
rect 210138 231192 211738 231592
rect 206938 229992 208538 230792
rect 206538 227592 208538 229992
rect 210138 228392 211338 231192
rect 214538 230792 216138 231592
rect 226938 231192 228538 231592
rect 228938 231192 230538 231592
rect 217338 230792 218538 231192
rect 214138 229992 215738 230792
rect 216938 230392 218538 230792
rect 216538 229992 218538 230392
rect 226938 230392 230538 231192
rect 231338 231592 232538 232392
rect 232938 231992 234538 232392
rect 246538 231592 250538 232792
rect 280938 232392 282938 233592
rect 283738 232392 286538 233592
rect 299738 233592 300538 233992
rect 301338 233592 302938 233992
rect 299738 233192 302938 233592
rect 299338 232792 303338 233192
rect 303738 232792 306938 233992
rect 310138 233592 311738 234392
rect 312938 233992 314538 234792
rect 312538 233592 314538 233992
rect 310138 233192 314938 233592
rect 299338 232392 302938 232792
rect 258138 231592 260938 231992
rect 272538 231592 275338 231992
rect 231338 230792 232938 231592
rect 246138 231192 250538 231592
rect 257738 231192 261738 231592
rect 271338 231192 276138 231592
rect 280938 231192 286538 232392
rect 299738 231992 302938 232392
rect 299338 231592 302938 231992
rect 246138 230792 250138 231192
rect 256538 230792 262938 231192
rect 270138 230792 277338 231192
rect 280938 230792 284138 231192
rect 230938 230392 232938 230792
rect 233738 230392 234538 230792
rect 246138 230392 250538 230792
rect 255338 230392 263738 230792
rect 269338 230392 277738 230792
rect 280938 230392 283738 230792
rect 284538 230392 286538 231192
rect 298938 230792 303338 231592
rect 305338 231192 306938 232792
rect 309338 232392 314938 233192
rect 308938 231992 314938 232392
rect 315738 233192 317338 234792
rect 320538 235192 321738 236792
rect 323338 235992 324938 237192
rect 323738 235592 324938 235992
rect 320538 234392 322138 235192
rect 323738 234792 325338 235592
rect 320938 233592 322138 234392
rect 308938 231592 314538 231992
rect 308938 231192 311338 231592
rect 312538 231192 314538 231592
rect 315738 231192 316938 233192
rect 320938 232792 322538 233592
rect 321338 231592 322538 232792
rect 324138 232792 325338 234792
rect 324138 231992 325738 232792
rect 298938 230392 300538 230792
rect 214138 229192 218938 229992
rect 226938 229592 228938 230392
rect 229338 229992 230138 230392
rect 230938 229592 234938 230392
rect 245738 229992 250538 230392
rect 254538 229992 264138 230392
rect 268538 229992 272938 230392
rect 274938 229992 278138 230392
rect 227338 229192 228938 229592
rect 214138 228792 217338 229192
rect 214538 228392 216538 228792
rect 217738 228392 218938 229192
rect 227738 228792 228938 229192
rect 231338 229192 234538 229592
rect 231338 228792 232538 229192
rect 232938 228792 234938 229192
rect 245338 228792 250538 229992
rect 253738 229592 257738 229992
rect 260938 229592 264938 229992
rect 267338 229592 271338 229992
rect 276138 229592 278538 229992
rect 253738 229192 256938 229592
rect 262138 229192 265338 229592
rect 267338 229192 270538 229592
rect 276938 229192 278538 229592
rect 253738 228792 256138 229192
rect 258538 228792 260538 229192
rect 262938 228792 265738 229192
rect 267338 228792 270138 229192
rect 272138 228792 274538 229192
rect 277338 228792 278938 229192
rect 280938 228792 283338 230392
rect 284538 229992 286138 230392
rect 284138 229192 285738 229992
rect 299338 229592 300538 230392
rect 298938 229192 300538 229592
rect 301338 229592 302938 230792
rect 303738 229992 306538 231192
rect 309338 230792 310138 231192
rect 312938 230792 314138 231192
rect 316138 230792 316938 231192
rect 317738 230792 318538 231192
rect 317338 230392 318938 230792
rect 227338 228392 228938 228792
rect 229738 228392 230938 228792
rect 231738 228392 232538 228792
rect 233338 228392 234938 228792
rect 245738 228392 249338 228792
rect 256938 228392 261338 228792
rect 263738 228392 265738 228792
rect 267738 228392 268938 228792
rect 270538 228392 276138 228792
rect 277738 228392 279338 228792
rect 209738 227592 211338 228392
rect 218138 227592 218938 228392
rect 226938 227592 228938 228392
rect 229338 227992 232538 228392
rect 232938 227992 235338 228392
rect 245738 227992 248138 228392
rect 256138 227992 261738 228392
rect 229338 227592 235338 227992
rect 246138 227592 247738 227992
rect 255738 227592 262538 227992
rect 264138 227592 265738 228392
rect 269738 227992 276538 228392
rect 278138 227992 279338 228392
rect 269338 227592 276938 227992
rect 278538 227592 279338 227992
rect 280938 228392 282938 228792
rect 283738 228392 285338 229192
rect 298938 228792 300938 229192
rect 301338 228792 302538 229592
rect 303738 229192 306938 229992
rect 280938 227592 285338 228392
rect 299338 228392 302538 228792
rect 299338 227992 302938 228392
rect 303338 227992 306938 229192
rect 316938 229592 318538 230392
rect 316938 229192 318138 229592
rect 316938 228792 317738 229192
rect 321738 228792 322938 231592
rect 324538 231192 325738 231992
rect 324538 228792 326138 231192
rect 322138 228392 322938 228792
rect 309338 227992 309738 228392
rect 313338 227992 313738 228392
rect 206538 215992 208138 227592
rect 210138 227192 210938 227592
rect 209738 224792 210938 227192
rect 216138 227192 219738 227592
rect 227338 227192 228538 227592
rect 216138 226392 222138 227192
rect 229738 226792 230538 227592
rect 230938 227192 232538 227592
rect 233338 227192 234938 227592
rect 246138 227192 248138 227592
rect 231338 226792 232938 227192
rect 233738 226792 234538 227192
rect 229738 226392 230938 226792
rect 231738 226392 232938 226792
rect 246538 226392 248138 227192
rect 254538 227192 262938 227592
rect 254538 226792 263338 227192
rect 250538 226392 251338 226792
rect 216538 225992 221738 226392
rect 227738 225992 229338 226392
rect 229738 225992 232938 226392
rect 216538 225592 220938 225992
rect 216538 224792 218538 225592
rect 209338 224392 210938 224792
rect 216138 224392 218538 224792
rect 209738 223192 210938 224392
rect 215738 223992 218538 224392
rect 215338 223192 218538 223992
rect 227738 225192 232938 225992
rect 246938 225192 248138 226392
rect 249738 225992 251338 226392
rect 254538 225992 260538 226792
rect 260938 225992 263738 226792
rect 249338 225192 251338 225992
rect 254938 225592 256538 225992
rect 256938 225592 263738 225992
rect 227738 224792 231338 225192
rect 232138 224792 232938 225192
rect 227738 223592 231738 224792
rect 233738 223592 235338 225192
rect 246538 223592 248138 225192
rect 248938 224792 251338 225192
rect 249338 223592 251338 224792
rect 255738 225192 256538 225592
rect 257338 225192 259338 225592
rect 259738 225192 263738 225592
rect 255738 224792 263738 225192
rect 255738 224392 263338 224792
rect 256138 223992 263338 224392
rect 256538 223592 263338 223992
rect 264538 223592 265738 227592
rect 268938 227192 277338 227592
rect 268538 226792 277738 227192
rect 280938 226792 285738 227592
rect 268138 226392 275338 226792
rect 268138 225192 270538 226392
rect 271338 225992 274538 226392
rect 275738 225992 277738 226792
rect 271338 225592 274138 225992
rect 274938 225592 277738 225992
rect 281338 226392 285738 226792
rect 298938 226392 300138 227992
rect 300938 227592 302938 227992
rect 300938 227192 303338 227592
rect 303738 227192 306538 227992
rect 301338 226792 306538 227192
rect 308938 227592 310138 227992
rect 308938 227192 310538 227592
rect 312538 227192 314138 227992
rect 308938 226792 310938 227192
rect 312138 226792 314138 227192
rect 301338 226392 302538 226792
rect 281338 225992 282938 226392
rect 283338 225992 285738 226392
rect 300938 225992 302538 226392
rect 271738 225192 273338 225592
rect 274538 225192 277338 225592
rect 268138 224792 270938 225192
rect 272138 224792 276938 225192
rect 268138 224392 276938 224792
rect 268538 223992 276938 224392
rect 269338 223592 276938 223992
rect 209338 222392 210938 223192
rect 214938 222392 216138 223192
rect 216538 222792 218538 223192
rect 219338 223192 220138 223592
rect 221738 223192 222538 223592
rect 228138 223192 231738 223592
rect 232938 223192 235338 223592
rect 219338 222792 220538 223192
rect 209738 221992 210938 222392
rect 214538 221992 216138 222392
rect 216938 222392 218538 222792
rect 218938 222392 220538 222792
rect 220938 222792 222938 223192
rect 220938 222392 223338 222792
rect 209738 221592 210538 221992
rect 209738 221192 210938 221592
rect 214538 221192 215738 221992
rect 216938 221592 223338 222392
rect 228138 221992 230138 223192
rect 230938 222792 231338 223192
rect 232538 222792 234538 223192
rect 246938 222792 248538 223592
rect 230938 222392 235738 222792
rect 247338 222392 248538 222792
rect 249738 223192 251338 223592
rect 256938 223192 262938 223592
rect 230538 221992 236138 222392
rect 247338 221992 248938 222392
rect 228138 221592 236538 221992
rect 247738 221592 248938 221992
rect 249738 221592 251738 223192
rect 258138 222792 259738 223192
rect 261338 222792 262938 223192
rect 260538 222392 262938 222792
rect 264138 222392 265738 223592
rect 270138 223192 276538 223592
rect 270938 222792 275738 223192
rect 271338 222392 274538 222792
rect 260138 221992 262538 222392
rect 259338 221592 262138 221992
rect 216938 221192 221738 221592
rect 209338 220392 210938 221192
rect 209738 219592 210938 220392
rect 209338 218792 210938 219592
rect 209738 215992 210938 218792
rect 214138 220392 215738 221192
rect 216538 220792 221738 221192
rect 216138 220392 221738 220792
rect 222138 220392 223738 221592
rect 228138 221192 236138 221592
rect 247738 221192 249338 221592
rect 214138 219192 221338 220392
rect 222538 219992 223738 220392
rect 214138 218392 216138 219192
rect 216938 218792 221738 219192
rect 222138 218792 223738 219992
rect 228538 220792 232138 221192
rect 233338 220792 236538 221192
rect 228538 219992 230538 220792
rect 231338 220392 232138 220792
rect 232938 220392 236538 220792
rect 248138 220792 249338 221192
rect 248138 220392 249738 220792
rect 230938 219992 236938 220392
rect 228538 219592 232938 219992
rect 233338 219592 236938 219992
rect 228938 219192 232938 219592
rect 233738 219192 236938 219592
rect 248538 219992 249738 220392
rect 250138 219992 251738 221592
rect 258938 221192 261338 221592
rect 258938 220792 260538 221192
rect 264138 220392 265338 222392
rect 272138 221992 275738 222392
rect 281338 221992 282538 225992
rect 283738 225592 285338 225992
rect 284138 223592 285338 225592
rect 300538 225192 302538 225992
rect 302938 225992 306538 226792
rect 308538 226392 311338 226792
rect 311738 226392 314538 226792
rect 302938 225192 306138 225992
rect 298538 224392 299738 225192
rect 300938 224792 303738 225192
rect 304138 224792 306138 225192
rect 283738 222392 285338 223592
rect 298138 223592 299738 224392
rect 300538 223992 302138 224792
rect 302538 223992 306138 224792
rect 308538 225592 314538 226392
rect 315738 226392 316938 228392
rect 315738 225992 317338 226392
rect 315338 225592 317338 225992
rect 308538 224792 317338 225592
rect 298138 223192 300138 223592
rect 300538 223192 305738 223992
rect 298538 222792 305738 223192
rect 299338 222392 301338 222792
rect 272538 221592 276138 221992
rect 281338 221592 282138 221992
rect 283738 221592 284938 222392
rect 297738 221992 298938 222392
rect 299738 221992 301338 222392
rect 301738 221992 303338 222792
rect 303738 221992 305338 222792
rect 273738 221192 274938 221592
rect 280938 220392 282138 221592
rect 283338 221192 284938 221592
rect 297338 221592 300938 221992
rect 301738 221592 305338 221992
rect 308538 222392 312138 224792
rect 312938 224392 317338 224792
rect 312938 223592 314938 224392
rect 312938 222792 314538 223592
rect 308538 221592 310138 222392
rect 310938 221992 312138 222392
rect 313338 221992 314538 222792
rect 315738 222792 317338 224392
rect 322138 225992 323338 228392
rect 322138 225192 323738 225992
rect 324938 225592 326538 228792
rect 322138 223992 323338 225192
rect 322138 223592 323738 223992
rect 322538 223192 323738 223592
rect 322538 222792 323338 223192
rect 313338 221592 314138 221992
rect 315738 221592 316938 222792
rect 322538 222392 323738 222792
rect 297338 221192 300538 221592
rect 301338 221192 302538 221592
rect 283338 220392 284538 221192
rect 297338 220792 300938 221192
rect 301338 220792 302138 221192
rect 296938 220392 298538 220792
rect 298938 220392 302138 220792
rect 302938 220392 304938 221592
rect 308938 221192 309738 221592
rect 280938 219992 281738 220392
rect 282938 219992 284538 220392
rect 296538 219992 298138 220392
rect 298938 219992 304538 220392
rect 248538 219192 251738 219992
rect 280538 219192 281738 219992
rect 282538 219192 284138 219992
rect 296538 219592 300538 219992
rect 300938 219592 304538 219992
rect 307338 219592 308938 219992
rect 296538 219192 300138 219592
rect 301338 219192 304538 219592
rect 306538 219192 312538 219592
rect 322138 219192 323738 222392
rect 228938 218792 231338 219192
rect 231738 218792 232538 219192
rect 216938 218392 223338 218792
rect 229338 218392 231338 218792
rect 214138 217992 215738 218392
rect 213738 217592 215338 217992
rect 217338 217592 223338 218392
rect 229738 217592 231338 218392
rect 232138 218392 233338 218792
rect 234138 218392 235738 219192
rect 232138 217992 235738 218392
rect 236538 217992 238138 218792
rect 248538 218392 252138 219192
rect 280138 218792 281338 219192
rect 282138 218792 283738 219192
rect 296538 218792 301738 219192
rect 232138 217592 235338 217992
rect 214138 217192 214938 217592
rect 217338 217192 220138 217592
rect 220938 217192 223338 217592
rect 230138 217192 235738 217592
rect 236538 217192 238538 217992
rect 248938 217592 252138 218392
rect 262938 218392 263738 218792
rect 262938 217992 264138 218392
rect 280138 217992 283338 218792
rect 296138 218392 297738 218792
rect 298138 218392 302138 218792
rect 302538 218392 304138 219192
rect 306138 218792 312938 219192
rect 305738 218392 312538 218792
rect 295738 217992 297338 218392
rect 298138 217992 303738 218392
rect 305738 217992 307338 218392
rect 307738 217992 312538 218392
rect 322138 217992 323338 219192
rect 325338 218792 326538 225592
rect 262538 217592 264138 217992
rect 249338 217192 252538 217592
rect 217338 216792 218138 217192
rect 219338 216792 220138 217192
rect 221338 216392 222538 217192
rect 230138 216792 234138 217192
rect 230538 216392 232538 216792
rect 232938 216392 234138 216792
rect 234538 216392 238538 217192
rect 249738 216792 252538 217192
rect 250938 216392 252538 216792
rect 262138 216792 263738 217592
rect 268938 217192 270138 217992
rect 279738 217592 282938 217992
rect 279738 217192 282538 217592
rect 295338 217192 297338 217992
rect 299738 217592 303738 217992
rect 300138 217192 303338 217592
rect 308138 217192 309738 217992
rect 316938 217592 317738 217992
rect 322138 217592 323738 217992
rect 312938 217192 314938 217592
rect 316138 217192 318538 217592
rect 268938 216792 270538 217192
rect 279738 216792 281738 217192
rect 295738 216792 296938 217192
rect 300938 216792 303338 217192
rect 262138 216392 264938 216792
rect 266938 216392 270538 216792
rect 220538 215992 222938 216392
rect 230538 215992 236938 216392
rect 237338 215992 238138 216392
rect 206538 214792 208538 215992
rect 209738 215192 211338 215992
rect 219738 215592 223338 215992
rect 230938 215592 236938 215992
rect 251338 215592 252938 216392
rect 262138 215992 270538 216392
rect 279338 216392 280938 216792
rect 299338 216392 303338 216792
rect 308538 216392 309738 217192
rect 312538 216792 318538 217192
rect 279338 215992 280538 216392
rect 262138 215592 270138 215992
rect 278938 215592 280538 215992
rect 296938 215592 298538 216392
rect 299338 215592 302938 216392
rect 219738 215192 221738 215592
rect 222138 215192 223738 215592
rect 206938 212392 208538 214792
rect 210138 212392 211338 215192
rect 219338 214792 221338 215192
rect 222538 214792 223738 215192
rect 230938 214792 234938 215592
rect 235738 215192 237338 215592
rect 238938 215192 240138 215592
rect 235738 214792 237738 215192
rect 238538 214792 240538 215192
rect 251738 214792 253338 215592
rect 262538 215192 267738 215592
rect 278938 215192 280138 215592
rect 265338 214792 266938 215192
rect 278538 214792 280138 215192
rect 293738 214792 295338 215592
rect 296538 215192 302938 215592
rect 308538 215992 310538 216392
rect 312138 215992 318938 216792
rect 308538 215592 311338 215992
rect 312138 215592 313738 215992
rect 308538 215192 311738 215592
rect 312138 215192 313338 215592
rect 218938 213992 220938 214792
rect 222938 214392 224138 214792
rect 223338 213992 223738 214392
rect 231338 213992 233338 214792
rect 233738 214392 237738 214792
rect 238138 214392 240538 214792
rect 234138 213992 240538 214392
rect 252138 214392 253338 214792
rect 252138 213992 253738 214392
rect 264938 213992 266138 214392
rect 266538 213992 266938 214392
rect 278538 213992 279738 214792
rect 293738 214392 295738 214792
rect 296538 214392 302538 215192
rect 308938 214792 313338 215192
rect 310138 214392 313338 214792
rect 293738 213992 297338 214392
rect 298538 213992 302538 214392
rect 308938 213992 311738 214392
rect 218938 213592 220538 213992
rect 207338 210392 208938 212392
rect 210138 211592 211738 212392
rect 207738 209192 208938 210392
rect 210538 210792 211738 211592
rect 218538 211192 220538 213592
rect 231738 213192 233738 213992
rect 234138 213592 236138 213992
rect 236538 213592 240938 213992
rect 252538 213592 254138 213992
rect 234538 213192 235738 213592
rect 236538 213192 238938 213592
rect 240138 213192 241338 213592
rect 252938 213192 254138 213592
rect 231738 212792 234138 213192
rect 222138 212392 222538 212792
rect 232138 212392 234138 212792
rect 236938 212792 238938 213192
rect 239738 212792 241738 213192
rect 252938 212792 254538 213192
rect 264938 212792 267338 213992
rect 278138 213592 279338 213992
rect 292538 213592 297338 213992
rect 299338 213592 302138 213992
rect 277738 212792 278938 213592
rect 292138 213192 294538 213592
rect 294938 213192 296938 213592
rect 291738 212792 296938 213192
rect 299738 213192 302138 213592
rect 308138 213592 311738 213992
rect 312138 213992 313338 214392
rect 314538 213992 316938 215992
rect 317738 215592 318938 215992
rect 322138 215192 323338 217592
rect 324938 215592 326538 218792
rect 322138 214792 322938 215192
rect 312138 213592 316938 213992
rect 308138 213192 311338 213592
rect 312538 213192 319338 213592
rect 299738 212792 301738 213192
rect 236938 212392 239338 212792
rect 239738 212392 242138 212792
rect 210538 209592 212138 210792
rect 218538 209992 220938 211192
rect 221738 210792 223338 212392
rect 232538 211992 234538 212392
rect 237338 211992 239338 212392
rect 240138 211992 242138 212392
rect 253338 212392 254538 212792
rect 263738 212392 266938 212792
rect 268538 212392 270538 212792
rect 253338 211992 254938 212392
rect 263338 211992 266538 212392
rect 267738 211992 270938 212392
rect 277338 211992 278538 212792
rect 291338 212392 297738 212792
rect 298938 212392 301738 212792
rect 307738 212792 310138 213192
rect 312938 212792 319338 213192
rect 307738 212392 309738 212792
rect 313338 212392 314938 212792
rect 315738 212392 319338 212792
rect 290938 211992 293338 212392
rect 294138 211992 296138 212392
rect 296538 211992 301338 212392
rect 232538 211592 234938 211992
rect 235738 211592 236938 211992
rect 237738 211592 239738 211992
rect 240538 211592 242938 211992
rect 232938 210792 237338 211592
rect 237738 211192 242938 211592
rect 253738 211592 254938 211992
rect 253738 211192 255338 211592
rect 261738 211192 270938 211992
rect 276938 211592 278138 211992
rect 290938 211592 292938 211992
rect 293738 211592 295738 211992
rect 296538 211592 300538 211992
rect 276938 211192 277738 211592
rect 290938 211192 295338 211592
rect 296138 211192 300538 211592
rect 238138 210792 243338 211192
rect 254138 210792 255738 211192
rect 261738 210792 270138 211192
rect 276538 210792 277738 211192
rect 291338 210792 294938 211192
rect 295738 210792 300138 211192
rect 221738 210392 225338 210792
rect 233338 210392 237338 210792
rect 238538 210392 243338 210792
rect 254538 210392 255738 210792
rect 267338 210392 269738 210792
rect 221338 209992 225738 210392
rect 233738 209992 238138 210392
rect 238938 209992 243738 210392
rect 254538 209992 256138 210392
rect 264938 209992 269338 210392
rect 276138 209992 277338 210792
rect 289338 210392 290938 210792
rect 292538 210392 296538 210792
rect 288938 209992 290938 210392
rect 292938 209992 296538 210392
rect 297338 210392 300138 210792
rect 297338 209992 299738 210392
rect 207738 207992 209338 209192
rect 210938 208792 212138 209592
rect 218938 209592 225738 209992
rect 234138 209592 236138 209992
rect 236538 209592 238538 209992
rect 238938 209592 240538 209992
rect 241738 209592 244138 209992
rect 254938 209592 256538 209992
rect 218938 209192 225338 209592
rect 234138 209192 238538 209592
rect 239738 209192 240138 209592
rect 242138 209192 244538 209592
rect 254938 209192 256938 209592
rect 219338 208792 225338 209192
rect 234538 208792 238538 209192
rect 241738 208792 246138 209192
rect 255338 208792 256938 209192
rect 264538 208792 268938 209992
rect 275738 209592 276938 209992
rect 275338 209192 276938 209592
rect 288938 209592 291338 209992
rect 294538 209592 296538 209992
rect 296938 209592 299338 209992
rect 288938 209192 292138 209592
rect 293738 209192 294938 209592
rect 296938 209192 298938 209592
rect 208138 206392 209738 207992
rect 211338 207192 212538 208792
rect 219738 208392 224938 208792
rect 234938 208392 238538 208792
rect 240938 208392 246538 208792
rect 255338 208392 257338 208792
rect 264138 208392 268938 208792
rect 274938 208792 276938 209192
rect 287738 208792 288538 209192
rect 289338 208792 292138 209192
rect 293338 208792 294938 209192
rect 296538 208792 298538 209192
rect 274938 208392 276538 208792
rect 287338 208392 288938 208792
rect 289738 208392 292138 208792
rect 220138 207992 224138 208392
rect 234938 207992 237338 208392
rect 238938 207992 239738 208392
rect 240538 207992 242938 208392
rect 220538 207592 223738 207992
rect 235338 207592 237338 207992
rect 238538 207592 242938 207992
rect 243738 207992 246538 208392
rect 255738 207992 257738 208392
rect 264138 207992 269338 208392
rect 274538 207992 276538 208392
rect 286938 207992 288938 208392
rect 290938 207992 291738 208392
rect 292938 207992 295338 208792
rect 296138 208392 298538 208792
rect 295738 207992 298138 208392
rect 307738 207992 309338 212392
rect 310138 211992 311338 212392
rect 316138 211992 318938 212392
rect 310138 211592 311738 211992
rect 309738 208792 311738 211592
rect 316538 211592 318938 211992
rect 321738 211592 322938 214792
rect 324538 213592 326538 215592
rect 324538 212392 326138 213592
rect 324138 211592 326138 212392
rect 316538 211192 318538 211592
rect 316538 210792 318138 211192
rect 321338 210792 322538 211592
rect 316138 209992 318138 210792
rect 316138 209592 318538 209992
rect 316538 209192 318538 209592
rect 320938 209592 322538 210792
rect 324138 209992 325738 211592
rect 324138 209592 325338 209992
rect 310138 208392 311338 208792
rect 316938 208392 318938 209192
rect 320938 208792 322138 209592
rect 243738 207592 247338 207992
rect 255738 207592 258138 207992
rect 266538 207592 269338 207992
rect 274138 207592 276538 207992
rect 285738 207592 288538 207992
rect 292138 207592 298138 207992
rect 220938 207192 222938 207592
rect 235338 207192 237738 207592
rect 238138 207192 242938 207592
rect 244138 207192 245338 207592
rect 246138 207192 247738 207592
rect 256138 207192 258538 207592
rect 273738 207192 276538 207592
rect 211338 206392 212938 207192
rect 220538 206792 222538 207192
rect 236138 206792 240138 207192
rect 240938 206792 243338 207192
rect 244938 206792 245738 207192
rect 246138 206792 248138 207192
rect 256138 206792 258938 207192
rect 273338 206792 276538 207192
rect 285338 206792 286938 207592
rect 287738 207192 288138 207592
rect 291738 207192 297738 207592
rect 287738 206792 288938 207192
rect 291738 206792 293738 207192
rect 294938 206792 297338 207192
rect 220538 206392 224138 206792
rect 236538 206392 239738 206792
rect 240538 206392 243738 206792
rect 208538 205192 210138 206392
rect 211738 205592 212938 206392
rect 220938 205992 224538 206392
rect 236538 205992 238938 206392
rect 240138 205992 243738 206392
rect 244938 205992 248538 206792
rect 256538 206392 259338 206792
rect 272938 206392 276538 206792
rect 285738 206392 286538 206792
rect 287338 206392 289338 206792
rect 290538 206392 293338 206792
rect 294538 206392 296938 206792
rect 248938 205992 250138 206392
rect 256538 205992 259738 206392
rect 272538 205992 276538 206392
rect 286938 205992 289338 206392
rect 221738 205592 224938 205992
rect 236938 205592 239338 205992
rect 240138 205592 244138 205992
rect 244938 205592 250938 205992
rect 256538 205592 260538 205992
rect 271738 205592 276538 205992
rect 283338 205592 284138 205992
rect 286138 205592 289338 205992
rect 208938 204792 210138 205192
rect 212138 204792 213338 205592
rect 222938 205192 224938 205592
rect 237338 205192 243738 205592
rect 245338 205192 250938 205592
rect 223338 204792 224938 205192
rect 237738 204792 241738 205192
rect 242538 204792 243338 205192
rect 245738 204792 246138 205192
rect 246938 204792 247738 205192
rect 248938 204792 250938 205192
rect 256938 205192 260938 205592
rect 270938 205192 276538 205592
rect 282938 205192 284538 205592
rect 285338 205192 289338 205592
rect 290138 205992 293338 206392
rect 294138 205992 296538 206392
rect 290138 205592 292138 205992
rect 293738 205592 296138 205992
rect 307338 205592 309338 207992
rect 317338 207192 318938 208392
rect 320538 207992 322138 208792
rect 323738 207992 325338 209592
rect 317338 206792 318538 207192
rect 316938 206392 318538 206792
rect 320538 206392 321738 207992
rect 323338 207592 325338 207992
rect 323338 206392 324938 207592
rect 316538 205992 318138 206392
rect 290138 205192 291738 205592
rect 293338 205192 295738 205592
rect 306938 205192 309338 205592
rect 316138 205592 317738 205992
rect 320138 205592 321338 206392
rect 316138 205192 317338 205592
rect 256938 204792 261338 205192
rect 270538 204792 276538 205192
rect 208938 203992 210538 204792
rect 212138 203992 213738 204792
rect 221338 204392 224938 204792
rect 220538 203992 224938 204392
rect 238138 203992 240938 204792
rect 242538 204392 243738 204792
rect 244938 204392 246138 204792
rect 248138 204392 248538 204792
rect 249738 204392 251738 204792
rect 256938 204392 262538 204792
rect 269338 204392 276538 204792
rect 280538 204392 281738 204792
rect 282538 204392 284138 205192
rect 284938 204792 287738 205192
rect 288538 204792 289738 205192
rect 290538 204792 291338 205192
rect 292938 204792 295338 205192
rect 305738 204792 308938 205192
rect 284938 204392 287338 204792
rect 288538 204392 290138 204792
rect 291738 204392 294938 204792
rect 304938 204392 308938 204792
rect 319738 204792 321338 205592
rect 322938 205992 324938 206392
rect 322938 204792 324538 205992
rect 319738 204392 320938 204792
rect 322938 204392 324138 204792
rect 242538 203992 244138 204392
rect 244538 203992 246538 204392
rect 247738 203992 248938 204392
rect 208938 203192 210938 203992
rect 209338 202792 210938 203192
rect 212538 203192 213738 203992
rect 220138 203592 224938 203992
rect 238538 203592 240938 203992
rect 242138 203592 246538 203992
rect 247338 203592 249338 203992
rect 250138 203592 252138 204392
rect 219738 203192 221738 203592
rect 222138 203192 224938 203592
rect 238938 203192 240938 203592
rect 241338 203192 249338 203592
rect 250538 203192 252138 203592
rect 256938 203992 263738 204392
rect 267738 203992 276938 204392
rect 256938 203592 276938 203992
rect 278138 203592 278938 203992
rect 279738 203592 281738 204392
rect 282938 203992 286538 204392
rect 286938 203992 290138 204392
rect 291338 203992 294538 204392
rect 304938 203992 308538 204392
rect 283338 203592 286138 203992
rect 286938 203592 289738 203992
rect 290938 203592 294138 203992
rect 304938 203592 306538 203992
rect 209338 201992 211338 202792
rect 212538 202392 214138 203192
rect 212938 201992 214138 202392
rect 219738 202392 220938 203192
rect 222538 202792 224938 203192
rect 229738 202792 231738 203192
rect 239338 202792 249338 203192
rect 249738 202792 253338 203192
rect 222538 202392 224538 202792
rect 229338 202392 232538 202792
rect 239738 202392 240138 202792
rect 240538 202392 250938 202792
rect 251738 202392 253338 202792
rect 254138 202392 255338 202792
rect 219738 201992 221338 202392
rect 222538 201992 224938 202392
rect 229738 201992 232538 202392
rect 240538 201992 248138 202392
rect 248938 201992 253338 202392
rect 209738 201192 211338 201992
rect 213338 201592 214538 201992
rect 219738 201592 225338 201992
rect 230938 201592 232938 201992
rect 210138 200392 211738 201192
rect 213338 200792 214938 201592
rect 220138 201192 225338 201592
rect 220538 200792 222138 201192
rect 223738 200792 225738 201192
rect 210138 199992 212138 200392
rect 210538 199592 212138 199992
rect 213738 199992 214938 200792
rect 224138 200392 226538 200792
rect 231738 200392 232938 201592
rect 240938 201592 247738 201992
rect 249338 201592 251738 201992
rect 252138 201592 253338 201992
rect 240938 201192 243338 201592
rect 244538 201192 247338 201592
rect 249338 201192 251338 201592
rect 252538 201192 253338 201592
rect 253738 201992 256538 202392
rect 256938 201992 259738 203592
rect 261338 203192 277338 203592
rect 277738 203192 279338 203592
rect 279738 203192 280938 203592
rect 281338 203192 282538 203592
rect 283338 203192 285338 203592
rect 286938 203192 288938 203592
rect 290138 203192 293338 203592
rect 261738 202792 279338 203192
rect 281338 202792 282938 203192
rect 283738 202792 285338 203192
rect 285738 202792 288538 203192
rect 289338 202792 292938 203192
rect 319338 202792 320538 204392
rect 322538 203192 324138 204392
rect 262538 202392 278938 202792
rect 280938 202392 283338 202792
rect 284138 202392 287738 202792
rect 288938 202392 292138 202792
rect 319338 202392 320138 202792
rect 263338 201992 278138 202392
rect 253738 201192 259738 201992
rect 263738 201592 278138 201992
rect 278538 201992 280538 202392
rect 281338 201992 283338 202392
rect 284938 201992 286938 202392
rect 288138 201992 291338 202392
rect 318938 201992 320138 202392
rect 322138 201992 323738 203192
rect 278538 201592 282938 201992
rect 283738 201592 284538 201992
rect 284938 201592 290938 201992
rect 318538 201592 320138 201992
rect 264538 201192 282138 201592
rect 283338 201192 290538 201592
rect 241338 200792 246938 201192
rect 241738 200392 246938 200792
rect 247738 200792 251338 201192
rect 252138 200792 259738 201192
rect 264938 200792 270938 201192
rect 272938 200792 276138 201192
rect 276538 200792 282138 201192
rect 247738 200392 249738 200792
rect 224938 199992 226938 200392
rect 231338 199992 232938 200392
rect 213738 199592 215338 199992
rect 225338 199592 228538 199992
rect 230938 199592 232938 199992
rect 242938 199992 246538 200392
rect 247338 199992 249738 200392
rect 242938 199592 245738 199992
rect 247738 199592 249738 199992
rect 250138 200392 255738 200792
rect 256138 200392 259738 200792
rect 265338 200392 270538 200792
rect 250138 199992 255338 200392
rect 256138 199992 257738 200392
rect 250138 199592 252938 199992
rect 210538 199192 212538 199592
rect 210938 198392 212538 199192
rect 214138 199192 215338 199592
rect 226138 199192 232538 199592
rect 242938 199192 246138 199592
rect 248138 199192 249738 199592
rect 250538 199192 253338 199592
rect 253738 199192 257738 199992
rect 214138 198792 215738 199192
rect 226538 198792 232538 199192
rect 243338 198792 246538 199192
rect 248938 198792 250138 199192
rect 250938 198792 257338 199192
rect 214538 198392 215738 198792
rect 227738 198392 231738 198792
rect 244138 198392 247738 198792
rect 210938 197992 212938 198392
rect 214538 197992 216138 198392
rect 228538 197992 231338 198392
rect 244538 197992 248538 198392
rect 249338 197992 251338 198792
rect 252538 198392 257338 198792
rect 252538 197992 256938 198392
rect 211338 197592 212938 197992
rect 211338 196792 213338 197592
rect 214938 197192 216138 197992
rect 244538 197592 248938 197992
rect 249738 197592 251738 197992
rect 252938 197592 256938 197992
rect 258138 197592 259738 200392
rect 265738 199992 269738 200392
rect 273338 199992 276138 200792
rect 276938 199992 279738 200792
rect 280138 199992 282138 200792
rect 282938 199992 285338 201192
rect 285738 200792 289338 201192
rect 318538 200792 319738 201592
rect 321738 201192 323338 201992
rect 321738 200792 322938 201192
rect 286138 200392 288938 200792
rect 286138 199992 288538 200392
rect 318138 199992 319338 200792
rect 321338 199992 322938 200792
rect 266138 199592 269338 199992
rect 266938 199192 268938 199592
rect 273738 198792 276138 199992
rect 277338 199192 283338 199992
rect 283738 199592 288138 199992
rect 317738 199592 319338 199992
rect 320938 199592 322938 199992
rect 283738 199192 287338 199592
rect 317738 199192 318938 199592
rect 277738 198792 282938 199192
rect 283738 198792 286938 199192
rect 317338 198792 318938 199192
rect 320938 198792 322538 199592
rect 274138 197992 276538 198792
rect 277738 198392 282538 198792
rect 283338 198392 286138 198792
rect 278138 197992 285338 198392
rect 317338 197992 318538 198792
rect 320538 197992 322138 198792
rect 246138 197192 251738 197592
rect 253738 197192 256538 197592
rect 215338 196792 251738 197192
rect 252138 196792 256538 197192
rect 257738 197192 259738 197592
rect 274538 197192 276938 197992
rect 278538 197592 284938 197992
rect 316938 197592 318538 197992
rect 278938 197192 284538 197592
rect 316938 197192 318138 197592
rect 320138 197192 321738 197992
rect 211738 195992 213738 196792
rect 215338 196392 256138 196792
rect 257738 196392 259338 197192
rect 274938 196392 277338 197192
rect 279338 196792 284938 197192
rect 285338 196792 285738 197192
rect 298138 196792 305338 197192
rect 314138 196792 317738 197192
rect 279738 196392 317738 196792
rect 319738 196792 321738 197192
rect 319738 196392 321338 196792
rect 215338 195992 255738 196392
rect 212138 195592 214138 195992
rect 212538 195192 214138 195592
rect 215738 195592 255738 195992
rect 257338 195592 259338 196392
rect 275338 195992 277738 196392
rect 280138 195992 317738 196392
rect 319338 195992 321338 196392
rect 275738 195592 278138 195992
rect 280938 195592 317338 195992
rect 319338 195592 320938 195992
rect 215738 195192 255338 195592
rect 212538 194392 214538 195192
rect 216138 194792 217738 195192
rect 216538 194392 217738 194792
rect 218938 194792 220938 195192
rect 221338 194792 225338 195192
rect 225738 194792 230138 195192
rect 212938 193592 214938 194392
rect 216538 193992 218138 194392
rect 218938 193992 220538 194792
rect 221338 193992 222938 194792
rect 223338 193992 227738 194792
rect 228138 194392 230138 194792
rect 230538 194392 232538 195192
rect 232938 194392 234938 195192
rect 228138 193992 229738 194392
rect 230538 193992 232138 194392
rect 232938 193992 234538 194392
rect 235338 193992 236938 195192
rect 237738 193992 239338 195192
rect 240138 193992 241738 195192
rect 242538 194392 246538 195192
rect 246938 194792 254938 195192
rect 256938 194792 258938 195592
rect 275738 195192 278938 195592
rect 280938 195192 316938 195592
rect 319338 195192 320538 195592
rect 276138 194792 294138 195192
rect 246938 194392 248938 194792
rect 249338 194392 254938 194792
rect 256538 194392 258538 194792
rect 242538 193992 244138 194392
rect 244938 193992 246538 194392
rect 247338 193992 248538 194392
rect 249338 193992 254538 194392
rect 256138 193992 258538 194392
rect 276538 194392 294138 194792
rect 276538 193992 292138 194392
rect 292538 193992 294138 194392
rect 294938 194792 298938 195192
rect 299338 194792 301338 195192
rect 294938 193992 296538 194792
rect 297338 193992 298938 194792
rect 299738 193992 301338 194792
rect 302138 193992 303738 195192
rect 304138 194392 306138 195192
rect 304538 193992 306138 194392
rect 306538 193992 308538 195192
rect 308938 194392 310938 195192
rect 311338 194392 313338 195192
rect 313738 194392 316938 195192
rect 318938 194792 320538 195192
rect 308938 193992 310538 194392
rect 311738 193992 312938 194392
rect 314138 193992 316538 194392
rect 318538 193992 320138 194792
rect 216938 193592 218138 193992
rect 249338 193592 284538 193992
rect 285738 193592 290538 193992
rect 213338 193192 215338 193592
rect 213738 192792 215338 193192
rect 217338 192792 218538 193592
rect 248538 193192 284938 193592
rect 286538 193192 291338 193592
rect 314538 193192 316138 193992
rect 318138 193192 319738 193992
rect 222138 192792 223738 193192
rect 226538 192792 227738 193192
rect 230538 192792 231738 193192
rect 234138 192792 235738 193192
rect 238538 192792 239738 193192
rect 242538 192792 243738 193192
rect 247738 192792 278538 193192
rect 278938 192792 285338 193192
rect 287338 192792 293738 193192
rect 296538 192792 297738 193192
rect 213738 192392 215738 192792
rect 217338 192392 218938 192792
rect 214138 191992 215738 192392
rect 217738 191992 219338 192392
rect 222138 191992 224138 192792
rect 226138 192392 228138 192792
rect 230138 192392 232138 192792
rect 225738 191992 228138 192392
rect 229738 191992 232138 192392
rect 214138 191592 216138 191992
rect 214538 191192 216538 191592
rect 218138 191192 219738 191992
rect 222138 191592 223738 191992
rect 226138 191592 228138 191992
rect 230138 191592 232138 191992
rect 234138 191592 236138 192792
rect 238138 191592 240138 192792
rect 242138 191592 244138 192792
rect 246538 192392 256938 192792
rect 275738 192392 285338 192792
rect 288538 192392 293738 192792
rect 296138 192392 297738 192792
rect 300138 192392 301738 193192
rect 304538 192792 305738 193192
rect 308538 192792 309738 193192
rect 304138 192392 306138 192792
rect 308138 192392 309738 192792
rect 312138 192792 313738 193192
rect 314538 192792 315738 193192
rect 245738 191992 258538 192392
rect 275738 191992 285738 192392
rect 289338 191992 294138 192392
rect 295738 191992 297738 192392
rect 299738 191992 302138 192392
rect 303738 191992 306138 192392
rect 307738 191992 310138 192392
rect 244938 191592 250138 191992
rect 251338 191592 260938 191992
rect 274938 191592 285738 191992
rect 290138 191592 294538 191992
rect 222538 191192 223338 191592
rect 226538 191192 227338 191592
rect 230538 191192 231738 191592
rect 234538 191192 235338 191592
rect 238538 191192 239738 191592
rect 242538 191192 248938 191592
rect 250938 191192 277338 191592
rect 277738 191192 279738 191592
rect 282138 191192 286538 191592
rect 286938 191192 289338 191592
rect 290938 191192 294938 191592
rect 296138 191192 297738 191992
rect 300138 191592 301738 191992
rect 303738 191592 305738 191992
rect 300138 191192 301338 191592
rect 304138 191192 305738 191592
rect 308138 191592 309738 191992
rect 312138 191592 315338 192792
rect 317738 192392 319338 193192
rect 317338 191992 318938 192392
rect 316938 191592 318938 191992
rect 308138 191192 309338 191592
rect 312138 191192 314938 191592
rect 316938 191192 318538 191592
rect 214938 190792 216538 191192
rect 218538 190792 219738 191192
rect 242138 190792 248138 191192
rect 250538 190792 279738 191192
rect 282538 190792 289738 191192
rect 291738 190792 295738 191192
rect 312538 190792 314538 191192
rect 316538 190792 318138 191192
rect 214938 190392 216938 190792
rect 218938 190392 220138 190792
rect 241738 190392 247338 190792
rect 250138 190392 252538 190792
rect 254138 190392 280138 190792
rect 282938 190392 284538 190792
rect 284938 190392 289738 190792
rect 292538 190392 296138 190792
rect 312938 190392 314138 190792
rect 215338 189592 217338 190392
rect 218938 189992 220538 190392
rect 224138 189992 225338 190392
rect 228138 189992 229338 190392
rect 232538 189992 233338 190392
rect 236138 189992 237338 190392
rect 240138 189992 245738 190392
rect 248938 189992 252938 190392
rect 257338 189992 280538 190392
rect 282938 189992 287738 190392
rect 215738 189192 217738 189592
rect 219338 189192 220938 189992
rect 216138 188792 217738 189192
rect 220138 188792 221338 189192
rect 223738 188792 225738 189992
rect 227738 188792 229738 189992
rect 232138 189592 233738 189992
rect 231738 188792 233738 189592
rect 235738 189592 237738 189992
rect 238938 189592 245338 189992
rect 246538 189592 253338 189992
rect 259738 189592 280938 189992
rect 282938 189592 286538 189992
rect 235738 189192 244138 189592
rect 245738 189192 253338 189592
rect 235738 188792 242538 189192
rect 243738 188792 250138 189192
rect 251738 188792 253338 189192
rect 216138 188392 218138 188792
rect 220138 188392 221738 188792
rect 224138 188392 225338 188792
rect 228138 188392 229338 188792
rect 232138 188392 233338 188792
rect 235738 188392 249338 188792
rect 216538 187992 218538 188392
rect 216938 187192 218938 187992
rect 220538 187592 222138 188392
rect 235738 187992 240938 188392
rect 242138 187992 249338 188392
rect 250138 187992 251338 188392
rect 252138 187992 253338 188792
rect 254138 189192 256538 189592
rect 264538 189192 270538 189592
rect 275738 189192 281738 189592
rect 282538 189192 286138 189592
rect 288138 189192 290138 190392
rect 292138 189992 292938 190392
rect 293338 189992 296938 190392
rect 298538 189992 299738 190392
rect 302538 189992 303738 190392
rect 306538 189992 307738 190392
rect 310938 189992 312138 190392
rect 312538 189992 314138 190392
rect 316138 190392 318138 190792
rect 316138 189992 317738 190392
rect 291738 189592 292938 189992
rect 294138 189592 297738 189992
rect 298138 189592 300138 189992
rect 302538 189592 304138 189992
rect 291738 189192 293338 189592
rect 294938 189192 300138 189592
rect 254138 188392 257338 189192
rect 258138 188792 260538 189192
rect 275738 188792 276938 189192
rect 277338 188792 286138 189192
rect 287338 188792 289738 189192
rect 257738 188392 260938 188792
rect 261738 188392 264138 188792
rect 265738 188392 267338 188792
rect 269738 188392 270938 188792
rect 272938 188392 274938 188792
rect 275338 188392 289338 188792
rect 254138 187992 254938 188392
rect 234538 187592 239738 187992
rect 241338 187592 246938 187992
rect 247738 187592 249338 187992
rect 249738 187592 253338 187992
rect 254538 187592 254938 187992
rect 256138 187992 264138 188392
rect 256138 187592 256938 187992
rect 257738 187592 258938 187992
rect 220938 187192 222538 187592
rect 226138 187192 227338 187592
rect 230138 187192 231338 187592
rect 233738 187192 238938 187592
rect 240538 187192 246138 187592
rect 217338 186792 219338 187192
rect 221338 186792 222938 187192
rect 217738 186392 219738 186792
rect 221738 186392 222938 186792
rect 218138 185992 220138 186392
rect 221738 185992 223738 186392
rect 226138 185992 227738 187192
rect 230138 186392 231738 187192
rect 232938 186792 238138 187192
rect 239738 186792 245338 187192
rect 247738 186792 253338 187592
rect 257738 187192 258538 187592
rect 259738 187192 262538 187992
rect 262938 187592 264138 187992
rect 260138 186792 260538 187192
rect 261338 186792 262138 187192
rect 263338 186792 264138 187592
rect 264938 187992 267738 188392
rect 268938 187992 271738 188392
rect 264938 187592 268138 187992
rect 268538 187592 271738 187992
rect 272538 187992 279738 188392
rect 280538 187992 289338 188392
rect 291338 187992 292938 189192
rect 295738 188792 300138 189192
rect 302138 188792 304138 189592
rect 306138 188792 308138 189992
rect 310538 189592 313738 189992
rect 315738 189592 317738 189992
rect 310138 189192 313338 189592
rect 315738 189192 317338 189592
rect 310538 188792 313338 189192
rect 315338 188792 316938 189192
rect 296138 188392 300138 188792
rect 302538 188392 303738 188792
rect 306538 188392 307738 188792
rect 310538 188392 312938 188792
rect 314938 188392 316938 188792
rect 296938 187992 300138 188392
rect 310938 187992 312538 188392
rect 314538 187992 316538 188392
rect 264938 187192 272138 187592
rect 272538 187192 275738 187992
rect 276138 187592 287738 187992
rect 291338 187592 293738 187992
rect 297738 187592 300538 187992
rect 310938 187592 312138 187992
rect 314538 187592 316138 187992
rect 276138 187192 287338 187592
rect 291738 187192 294138 187592
rect 298138 187192 300938 187592
rect 304538 187192 306138 187592
rect 308538 187192 309738 187592
rect 310538 187192 312138 187592
rect 314138 187192 315738 187592
rect 264938 186792 265738 187192
rect 266938 186792 268138 187192
rect 268538 186792 269738 187192
rect 270538 186792 271738 187192
rect 272538 186792 273338 187192
rect 274538 186792 275738 187192
rect 276538 186792 278138 187192
rect 278538 186792 282938 187192
rect 283338 186792 286938 187192
rect 292538 186792 294538 187192
rect 298538 186792 301338 187192
rect 232138 186392 236938 186792
rect 238938 186392 241338 186792
rect 242138 186392 244538 186792
rect 247738 186392 249338 186792
rect 252138 186392 253338 186792
rect 265338 186392 265738 186792
rect 267338 186392 267738 186792
rect 268938 186392 269338 186792
rect 270938 186392 271338 186792
rect 272538 186392 272938 186792
rect 274938 186392 275338 186792
rect 276938 186392 284538 186792
rect 230138 185992 236138 186392
rect 238138 185992 240938 186392
rect 242138 185992 244138 186392
rect 247738 185992 249738 186392
rect 251738 185992 255738 186392
rect 218138 185592 220538 185992
rect 218538 185192 220538 185592
rect 222538 185192 224138 185992
rect 226538 185592 227338 185992
rect 230538 185592 235338 185992
rect 237738 185592 240138 185992
rect 241338 185592 243738 185992
rect 247738 185592 256538 185992
rect 277338 185592 284538 186392
rect 285338 186392 286938 186792
rect 293338 186392 294538 186792
rect 297338 186392 298138 186792
rect 299338 186392 301738 186792
rect 285338 185592 287338 186392
rect 288938 185992 290538 186392
rect 288538 185592 290938 185992
rect 291738 185592 292938 185992
rect 293338 185592 294938 186392
rect 296938 185992 298938 186392
rect 299738 185992 302538 186392
rect 304138 185992 306138 187192
rect 308138 186792 312138 187192
rect 313738 186792 315738 187192
rect 308138 186392 311338 186792
rect 313338 186392 315338 186792
rect 296538 185592 299338 185992
rect 300538 185592 302938 185992
rect 304538 185592 305738 185992
rect 308538 185592 310938 186392
rect 313338 185992 314938 186392
rect 312938 185592 314938 185992
rect 230538 185192 234538 185592
rect 236538 185192 238938 185592
rect 240938 185192 243338 185592
rect 246938 185192 256538 185592
rect 257738 185192 260138 185592
rect 262138 185192 263738 185592
rect 266538 185192 267338 185592
rect 270538 185192 270938 185592
rect 273738 185192 275738 185592
rect 276938 185192 282538 185592
rect 283338 185192 284138 185592
rect 285738 185192 287338 185592
rect 218938 184792 220938 185192
rect 222938 184792 224538 185192
rect 230138 184792 234138 185192
rect 236138 184792 238138 185192
rect 240538 184792 242538 185192
rect 246538 184792 256538 185192
rect 219338 184392 221338 184792
rect 223338 184392 224938 184792
rect 229338 184392 233338 184792
rect 236138 184392 237338 184792
rect 239738 184392 242138 184792
rect 244138 184392 244938 184792
rect 246538 184392 252938 184792
rect 254138 184392 256138 184792
rect 257338 184392 260538 185192
rect 261338 184792 264138 185192
rect 265738 184792 268138 185192
rect 269738 184792 272138 185192
rect 273338 184792 276138 185192
rect 219738 183992 221738 184392
rect 223738 183992 225338 184392
rect 228938 183992 232538 184392
rect 238938 183992 241738 184392
rect 243738 183992 244938 184392
rect 219738 183592 222138 183992
rect 220138 183192 222138 183592
rect 224138 183592 225338 183992
rect 228538 183592 232138 183992
rect 237738 183592 241338 183992
rect 242938 183592 244938 183992
rect 246138 183992 248138 184392
rect 248538 183992 252938 184392
rect 257738 183992 260138 184392
rect 261338 183992 264538 184792
rect 265338 183992 268538 184792
rect 269338 184392 272538 184792
rect 269338 183992 272138 184392
rect 272938 183992 276138 184792
rect 276538 184792 281738 185192
rect 282938 184792 284538 185192
rect 288138 184792 291338 185592
rect 291738 185192 294938 185592
rect 298138 185192 299338 185592
rect 300938 185192 303338 185592
rect 308938 185192 310538 185592
rect 312538 185192 314538 185592
rect 292138 184792 294538 185192
rect 276538 184392 280138 184792
rect 276938 183992 280138 184392
rect 282938 184392 284938 184792
rect 290138 184392 291738 184792
rect 292538 184392 294138 184792
rect 298138 184392 299738 185192
rect 301338 184792 303738 185192
rect 308538 184792 310138 185192
rect 312538 184792 314138 185192
rect 302138 184392 304138 184792
rect 282938 183992 285338 184392
rect 289738 183992 291738 184392
rect 295338 183992 296138 184392
rect 297738 183992 299738 184392
rect 302538 183992 304938 184392
rect 308138 183992 309738 184792
rect 312138 184392 313738 184792
rect 311738 183992 313338 184392
rect 246138 183592 247738 183992
rect 224138 183192 225738 183592
rect 228138 183192 231338 183592
rect 236938 183192 240538 183592
rect 242538 183192 244938 183592
rect 245738 183192 247338 183592
rect 248538 183192 253338 183992
rect 258938 183592 259338 183992
rect 261738 183592 264138 183992
rect 265738 183592 268138 183992
rect 269738 183592 271738 183992
rect 273338 183592 275738 183992
rect 278138 183592 280138 183992
rect 266538 183192 267338 183592
rect 270538 183192 270938 183592
rect 274138 183192 275338 183592
rect 220538 182792 222538 183192
rect 220938 182392 222938 182792
rect 224938 182392 226538 183192
rect 227738 182792 230538 183192
rect 235338 182792 240138 183192
rect 241738 182792 244938 183192
rect 226938 182392 230138 182792
rect 233738 182392 239738 182792
rect 241338 182392 244938 182792
rect 245338 182792 247338 183192
rect 248138 182792 253338 183192
rect 259738 182792 260938 183192
rect 245338 182392 246938 182792
rect 247738 182392 253738 182792
rect 221338 181992 223338 182392
rect 225338 181992 229738 182392
rect 232938 181992 239338 182392
rect 240938 181992 246538 182392
rect 247738 181992 254138 182392
rect 221738 181592 223738 181992
rect 226138 181592 228938 181992
rect 231338 181592 234938 181992
rect 236538 181592 238938 181992
rect 240138 181592 242538 181992
rect 222138 181192 224138 181592
rect 226138 181192 228538 181592
rect 231338 181192 234138 181592
rect 236138 181192 238138 181592
rect 239738 181192 242138 181592
rect 222138 180792 224538 181192
rect 226538 180792 228138 181192
rect 231338 180792 233738 181192
rect 235738 180792 237738 181192
rect 239338 180792 241738 181192
rect 242938 180792 244538 181992
rect 244938 180792 246138 181992
rect 247338 181592 254138 181992
rect 259338 181992 261338 182792
rect 273738 181992 275738 183192
rect 247338 181192 254538 181592
rect 222538 180392 224938 180792
rect 227338 180392 228938 180792
rect 231738 180392 233738 180792
rect 234938 180392 237338 180792
rect 238938 180392 240938 180792
rect 242538 180392 245738 180792
rect 246938 180392 250938 181192
rect 222938 179992 225338 180392
rect 223338 179592 225738 179992
rect 227738 179592 229338 180392
rect 232138 179992 236938 180392
rect 238538 179992 240538 180392
rect 232538 179592 236138 179992
rect 238138 179592 240138 179992
rect 242538 179592 243738 180392
rect 244538 179592 245338 180392
rect 246538 179592 248538 180392
rect 223738 179192 226138 179592
rect 228538 179192 230538 179592
rect 232938 179192 235338 179592
rect 237738 179192 239738 179592
rect 242138 179192 243738 179592
rect 246138 179192 248538 179592
rect 248938 179592 250938 180392
rect 251338 180392 254538 181192
rect 259338 180792 261738 181992
rect 273338 181192 275738 181992
rect 272138 180792 277338 181192
rect 224138 178792 226538 179192
rect 228938 178792 230538 179192
rect 233338 178792 234538 179192
rect 237338 178792 239338 179192
rect 241738 178792 243338 179192
rect 246138 178792 248138 179192
rect 224538 178392 226938 178792
rect 229338 178392 230938 178792
rect 236938 178392 238938 178792
rect 241338 178392 243338 178792
rect 224938 177992 227338 178392
rect 230138 177992 231738 178392
rect 236538 177992 238538 178392
rect 241338 177992 242938 178392
rect 245738 177992 247738 178792
rect 248938 177992 250538 179592
rect 225338 177592 227738 177992
rect 225738 177192 228138 177592
rect 230538 177192 232138 177992
rect 236138 177192 238538 177992
rect 240938 177592 242538 177992
rect 240538 177192 242538 177592
rect 245338 177192 247338 177992
rect 248538 177192 250538 177992
rect 251338 179192 254938 180392
rect 258138 179992 262938 180792
rect 272138 180392 275738 180792
rect 271738 179992 275738 180392
rect 276138 179992 277338 180792
rect 278538 179992 280138 183592
rect 283738 182792 285338 183992
rect 287738 183592 291338 183992
rect 292538 183592 292938 183992
rect 286938 183192 291338 183592
rect 291738 183192 293738 183592
rect 294938 183192 296938 183992
rect 297738 183192 299338 183992
rect 302938 183592 305338 183992
rect 307338 183592 308938 183992
rect 311338 183592 313338 183992
rect 286138 182792 290538 183192
rect 290938 182792 294538 183192
rect 283338 182392 284938 182792
rect 282938 181992 284938 182392
rect 285738 182392 290138 182792
rect 290938 182392 294938 182792
rect 285738 181992 287738 182392
rect 288538 181992 288938 182392
rect 290938 181992 292538 182392
rect 293338 181992 295338 182392
rect 295738 181992 297338 183192
rect 297738 182792 298938 183192
rect 300138 182792 301338 183592
rect 303338 183192 305738 183592
rect 306938 183192 308538 183592
rect 310938 183192 312938 183592
rect 303738 182792 308538 183192
rect 310538 182792 312538 183192
rect 297738 181992 301338 182792
rect 304138 182392 308138 182792
rect 310138 182392 312138 182792
rect 304538 181992 307338 182392
rect 310138 181992 311738 182392
rect 282138 181592 284538 181992
rect 281738 181192 284138 181592
rect 285738 181192 287338 181992
rect 291338 181592 292538 181992
rect 293738 181592 297338 181992
rect 298138 181592 300938 181992
rect 304938 181592 307338 181992
rect 309338 181592 311338 181992
rect 294138 181192 297338 181592
rect 298538 181192 300538 181592
rect 304938 181192 306938 181592
rect 308938 181192 310938 181592
rect 281738 180792 283738 181192
rect 285738 180792 287738 181192
rect 294138 180792 297738 181192
rect 298938 180792 299338 181192
rect 304538 180792 306538 181192
rect 308538 180792 310538 181192
rect 258138 179592 261338 179992
rect 256938 179192 259338 179592
rect 259738 179192 261338 179592
rect 261738 179592 262938 179992
rect 271338 179592 273338 179992
rect 273738 179592 275338 179992
rect 251338 178392 255338 179192
rect 256538 178792 259338 179192
rect 256938 178392 258938 178792
rect 260138 178392 260938 179192
rect 261738 178392 264138 179592
rect 270938 179192 273338 179592
rect 270938 178792 272938 179192
rect 274138 178792 275338 179592
rect 276138 178792 280138 179992
rect 281338 179592 283338 180792
rect 284538 180392 284938 180792
rect 286538 180392 287738 180792
rect 291338 180392 300138 180792
rect 284138 179992 285338 180392
rect 289338 179992 302138 180392
rect 304138 179992 305738 180792
rect 308138 180392 310138 180792
rect 307738 179992 309738 180392
rect 283738 179592 285338 179992
rect 288538 179592 305338 179992
rect 307338 179592 309738 179992
rect 281738 179192 285338 179592
rect 287338 179192 294138 179592
rect 294538 179192 296538 179592
rect 297738 179192 304538 179592
rect 306938 179192 308938 179592
rect 271338 178392 271738 178792
rect 273738 178392 275738 178792
rect 251338 177992 256540 178392
rect 259338 177994 261338 178392
rect 259338 177992 261738 177994
rect 263338 177992 265738 178392
rect 268938 177992 272138 178392
rect 273338 177992 276138 178392
rect 276938 177992 280138 178792
rect 282138 178792 284938 179192
rect 286538 178792 292538 179192
rect 294538 178792 296938 179192
rect 299338 178792 304538 179192
rect 306538 178792 308538 179192
rect 282138 178392 284538 178792
rect 286138 178392 291738 178792
rect 294538 178392 297338 178792
rect 299738 178392 300938 178792
rect 301738 178392 304138 178792
rect 306138 178392 308538 178792
rect 285338 177992 288938 178392
rect 289738 177992 292538 178392
rect 294138 177992 297338 178392
rect 298938 177992 300938 178392
rect 301338 177992 303338 178392
rect 305738 177992 307738 178392
rect 226538 176792 228538 177192
rect 231338 176792 233338 177192
rect 236538 176792 239338 177192
rect 240538 176792 242138 177192
rect 245338 176792 246938 177192
rect 226938 176392 228938 176792
rect 231738 176392 233738 176792
rect 236938 176392 242138 176792
rect 244938 176392 246938 176792
rect 227338 175992 229338 176392
rect 232138 175992 234138 176392
rect 237338 175992 241738 176392
rect 227738 175592 230138 175992
rect 232938 175592 234938 175992
rect 238138 175592 241738 175992
rect 244938 175592 246538 176392
rect 228138 175192 230538 175592
rect 233338 175192 235338 175592
rect 238538 175192 241338 175592
rect 228538 174792 230938 175192
rect 233738 174792 236138 175192
rect 239338 174792 241338 175192
rect 244938 174792 246138 175592
rect 248538 175192 250138 177192
rect 251338 176792 253338 177992
rect 253738 177592 258138 177992
rect 258938 177592 261738 177992
rect 262938 177592 266138 177992
rect 268538 177592 272538 177992
rect 272938 177592 276138 177992
rect 253738 176792 261738 177592
rect 262538 177192 266538 177592
rect 262138 176792 266538 177192
rect 268538 177192 274538 177592
rect 274938 177192 276138 177592
rect 268538 176792 272538 177192
rect 272938 176792 276138 177192
rect 276538 176792 280138 177992
rect 284938 177592 288138 177992
rect 289738 177592 292938 177992
rect 284138 177192 287338 177592
rect 283738 176792 287338 177192
rect 289338 177192 292938 177592
rect 294138 177592 297738 177992
rect 298938 177592 302938 177992
rect 305338 177592 307338 177992
rect 294138 177192 295338 177592
rect 289338 176792 291338 177192
rect 229338 174392 231738 174792
rect 234538 174392 236538 174792
rect 240138 174392 240938 174792
rect 229738 173992 232138 174392
rect 234938 173992 237338 174392
rect 244538 173992 245738 174792
rect 248538 174392 249738 175192
rect 230138 173592 232538 173992
rect 235738 173592 237738 173992
rect 230538 173192 233338 173592
rect 236538 173192 238938 173592
rect 244538 173192 245338 173992
rect 248938 173192 249738 174392
rect 231338 172792 233738 173192
rect 236938 172792 239338 173192
rect 249338 172792 249738 173192
rect 231738 172392 234138 172792
rect 237738 172392 239738 172792
rect 251738 172392 253338 176792
rect 254138 176392 258538 176792
rect 254138 175992 258138 176392
rect 259338 175992 261738 176792
rect 262538 176392 266538 176792
rect 268938 176392 272138 176792
rect 273338 176392 275738 176792
rect 276938 176392 280138 176792
rect 282938 176392 288138 176792
rect 289338 176392 290938 176792
rect 291738 176392 295338 177192
rect 296138 177192 297738 177592
rect 298538 177192 302538 177592
rect 304938 177192 306938 177592
rect 296138 176792 301738 177192
rect 304538 176792 306538 177192
rect 296538 176392 301338 176792
rect 304138 176392 306138 176792
rect 262938 175992 266138 176392
rect 269738 175992 270938 176392
rect 273738 175992 275338 176392
rect 278138 175992 280138 176392
rect 282538 175992 288538 176392
rect 289338 175992 291338 176392
rect 291738 175992 294938 176392
rect 296538 175992 300938 176392
rect 303738 175992 305738 176392
rect 254138 175592 256138 175992
rect 254538 173592 256138 175592
rect 256938 175192 258938 175592
rect 260538 175192 260938 175992
rect 271338 175592 273338 175992
rect 262138 175192 264138 175592
rect 256938 174392 259338 175192
rect 260138 174792 260938 175192
rect 259738 174392 261338 174792
rect 257738 173992 261338 174392
rect 261738 174392 264138 175192
rect 270938 174792 273338 175592
rect 274538 175192 274938 175592
rect 266538 174392 267338 174792
rect 261738 173992 263338 174392
rect 266138 173992 267738 174392
rect 272138 173992 273338 174792
rect 254938 172392 256138 173592
rect 258138 173192 262938 173992
rect 265738 173592 267738 173992
rect 272538 173592 273338 173992
rect 273738 174792 275338 175192
rect 276138 174792 280138 175992
rect 282138 175592 284538 175992
rect 285338 175592 288938 175992
rect 289338 175592 290938 175992
rect 292138 175592 294938 175992
rect 281738 175192 284138 175592
rect 285338 175192 290938 175592
rect 292538 175192 294538 175592
rect 296938 175192 300138 175992
rect 302938 175592 305338 175992
rect 302538 175192 304938 175592
rect 281338 174792 283738 175192
rect 273738 174392 275738 174792
rect 276138 174392 277338 174792
rect 273738 173992 277338 174392
rect 278538 174392 280138 174792
rect 280938 174392 282938 174792
rect 285338 174392 286938 175192
rect 287738 174792 290938 175192
rect 292938 174792 294138 175192
rect 294938 174792 299338 175192
rect 301738 174792 304538 175192
rect 288138 174392 290538 174792
rect 292538 174392 298538 174792
rect 301338 174392 303738 174792
rect 278538 173992 282938 174392
rect 285738 173992 286938 174392
rect 288538 173992 290138 174392
rect 291338 173992 298138 174392
rect 300938 173992 303338 174392
rect 273738 173592 276938 173992
rect 278538 173592 284138 173992
rect 285738 173592 287338 173992
rect 290538 173592 297338 173992
rect 300138 173592 302938 173992
rect 232538 171992 234938 172392
rect 238138 171992 240938 172392
rect 232938 171592 235738 171992
rect 238938 171592 241338 171992
rect 233338 171192 236138 171592
rect 239738 171192 242538 171592
rect 234138 170792 236938 171192
rect 240538 170792 243338 171192
rect 252138 170792 252938 172392
rect 254938 171992 256538 172392
rect 255338 171192 256138 171992
rect 259338 171592 261738 173192
rect 265738 172792 268138 173592
rect 265738 172392 268538 172792
rect 273738 172392 276138 173592
rect 278538 172792 287338 173592
rect 289338 173192 296938 173592
rect 299738 173192 302538 173592
rect 288538 172792 296138 173192
rect 298938 172792 302138 173192
rect 278138 172392 281338 172792
rect 281738 172392 287338 172792
rect 288138 172392 292138 172792
rect 292938 172392 295738 172792
rect 298538 172392 301338 172792
rect 264938 171992 265338 172392
rect 265738 171992 269338 172392
rect 264538 171592 269338 171992
rect 273738 171592 275738 172392
rect 278138 171992 280938 172392
rect 282138 171992 283338 172392
rect 284538 171992 290938 172392
rect 292538 171992 294138 172392
rect 297738 171992 300938 172392
rect 278138 171592 280538 171992
rect 282138 171592 283738 171992
rect 284938 171592 290138 171992
rect 291338 171592 294138 171992
rect 296938 171592 300138 171992
rect 259338 171192 261338 171592
rect 260138 170792 261338 171192
rect 264538 171192 269738 171592
rect 274138 171192 275338 171592
rect 278138 171192 280138 171592
rect 282138 171192 284138 171592
rect 286538 171192 289738 171592
rect 290938 171192 293738 171592
rect 296538 171192 299738 171592
rect 264538 170792 265738 171192
rect 266138 170792 267738 171192
rect 234938 170392 237738 170792
rect 241338 170392 244138 170792
rect 235338 169992 238138 170392
rect 242138 169992 244938 170392
rect 252138 169992 252538 170792
rect 263738 170392 265738 170792
rect 263338 169992 265738 170392
rect 266538 170392 267738 170792
rect 268138 170792 269738 171192
rect 277738 170792 280138 171192
rect 268138 170392 270538 170792
rect 266538 169992 267338 170392
rect 268538 169992 270938 170392
rect 277738 169992 279738 170792
rect 280938 169992 281738 170392
rect 282538 169992 284538 171192
rect 285738 170792 288938 171192
rect 289338 170792 292538 171192
rect 295738 170792 298938 171192
rect 285338 170392 292138 170792
rect 294938 170392 298538 170792
rect 284938 169992 290938 170392
rect 294538 169992 297738 170392
rect 236138 169592 239338 169992
rect 242938 169592 246138 169992
rect 263738 169592 264938 169992
rect 266138 169592 267738 169992
rect 268938 169592 270538 169992
rect 277338 169592 279338 169992
rect 280138 169592 290138 169992
rect 293738 169592 297338 169992
rect 236938 169192 239738 169592
rect 243338 169192 247338 169592
rect 261738 169192 264538 169592
rect 237338 168792 240538 169192
rect 244938 168792 248138 169192
rect 261338 168792 264538 169192
rect 265738 169192 268138 169592
rect 269738 169192 272538 169592
rect 277338 169192 289338 169592
rect 292938 169192 296538 169592
rect 265738 168792 268538 169192
rect 269338 168792 272938 169192
rect 277338 168792 288538 169192
rect 292138 168792 295738 169192
rect 238138 168392 241738 168792
rect 246138 168392 249738 168792
rect 260538 168392 266538 168792
rect 266938 168392 268538 168792
rect 238938 167992 242538 168392
rect 246538 167992 250938 168392
rect 260938 167992 268538 168392
rect 268938 167992 273338 168792
rect 239738 167592 243338 167992
rect 248138 167592 251738 167992
rect 252138 167592 252538 167992
rect 260938 167592 264938 167992
rect 240938 167192 244138 167592
rect 249738 167192 254538 167592
rect 261338 167192 264138 167592
rect 265738 167192 268138 167992
rect 268938 167592 272938 167992
rect 276938 167592 278538 168792
rect 279338 168392 280538 168792
rect 282538 168392 287338 168792
rect 291338 168392 294938 168792
rect 279738 167992 280138 168392
rect 282138 167992 286538 168392
rect 290538 167992 294538 168392
rect 280538 167592 285338 167992
rect 289738 167592 293738 167992
rect 269738 167192 272538 167592
rect 276938 167192 278138 167592
rect 278938 167192 283738 167592
rect 288538 167192 292538 167592
rect 241338 166792 245338 167192
rect 250138 166792 256138 167192
rect 266538 166792 267338 167192
rect 276538 166792 282138 167192
rect 287338 166792 292138 167192
rect 242538 166392 246138 166792
rect 251738 166392 256938 166792
rect 275338 166392 281338 166792
rect 286538 166392 290938 166792
rect 243738 165992 247338 166392
rect 253338 165992 261738 166392
rect 270138 165992 270938 166392
rect 271738 165992 279738 166392
rect 284938 165992 290138 166392
rect 244538 165592 248538 165992
rect 255338 165592 278138 165992
rect 283738 165592 289338 165992
rect 245338 165192 249738 165592
rect 256938 165192 276538 165592
rect 282938 165192 288538 165592
rect 246938 164792 251338 165192
rect 260938 164792 261738 165192
rect 262138 164792 271338 165192
rect 271738 164792 272538 165192
rect 280938 164792 286938 165192
rect 247738 164392 252938 164792
rect 266538 164392 266938 164792
rect 279338 164392 286138 164792
rect 248938 163992 254138 164392
rect 278138 163992 284938 164392
rect 250938 163592 256538 163992
rect 274938 163592 283338 163992
rect 251738 163192 259738 163592
rect 271338 163192 282138 163592
rect 253338 162792 262538 163192
rect 266138 162792 280538 163192
rect 255738 162392 277738 162792
rect 257338 161992 276138 162392
rect 260538 161592 273338 161992
rect 196984 151884 218276 157884
rect 196984 146172 202984 151884
rect 212276 146172 218276 151884
rect 196984 140172 218276 146172
rect 196984 129616 202984 140172
rect 212276 129616 218276 140172
rect 221222 135512 227222 157780
rect 236514 135512 242514 157780
rect 245282 151884 266574 157882
rect 221222 129512 242514 135512
rect 252717 129151 258715 151884
rect 269140 147836 275140 158104
rect 284432 147836 290432 158104
rect 294502 151906 315428 157906
rect 318502 151906 339428 157906
rect 309428 147964 315428 151906
rect 333428 147964 339428 151906
rect 269140 141836 290432 147836
rect 269140 129836 275138 141836
rect 284432 129836 290432 141836
rect 294912 141964 315428 147964
rect 318912 141964 339428 147964
rect 294912 136006 300912 141964
rect 318912 136006 324912 141964
rect 294912 130006 315568 136006
rect 318912 130006 339568 136006
<< fillblock >>
rect 165394 553901 200396 570901
rect 138394 512901 200396 553901
rect 415918 517730 517918 598730
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use LDO  LDO_0
timestamp 1667842615
transform -1 0 550078 0 -1 694876
box -8958 -8682 15320 8530
use decoupling_cell  decoupling_cell_0
timestamp 1668785275
transform 1 0 368582 0 1 242038
box 0 0 201600 203879
use mirrors  mirrors_0
timestamp 1668275587
transform 0 -1 358618 1 0 616664
box -18962 22 70826 31618
use pwm_lower  pwm_lower_0
timestamp 1668298669
transform 0 1 413660 -1 0 697163
box 4398 -2478 18637 19086
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_0
timestamp 1667857442
transform 1 0 335699 0 1 389400
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_1
timestamp 1667857442
transform 1 0 334699 0 1 389400
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_2
timestamp 1667857442
transform 1 0 468123 0 1 450054
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_3
timestamp 1667857442
transform 1 0 469123 0 1 450054
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_4
timestamp 1667857442
transform 1 0 54011 0 1 145689
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_5
timestamp 1667857442
transform 1 0 55011 0 1 145689
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_6
timestamp 1667857442
transform 1 0 56011 0 1 145689
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_7
timestamp 1667857442
transform 1 0 57011 0 1 145689
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_8
timestamp 1667857442
transform 1 0 60759 0 1 145778
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_9
timestamp 1667857442
transform 1 0 61759 0 1 145778
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_10
timestamp 1667857442
transform 1 0 62759 0 1 145778
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_11
timestamp 1667857442
transform 1 0 63759 0 1 145778
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_12
timestamp 1667857442
transform 1 0 551758 0 1 146748
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_13
timestamp 1667857442
transform 1 0 552758 0 1 146748
box -423 -423 423 423
use sky130_fd_pr__nfet_01v8_CY273Z  sky130_fd_pr__nfet_01v8_CY273Z_0
timestamp 1668290293
transform 0 1 57970 -1 0 147676
box -496 -260 496 260
use sky130_fd_pr__nfet_01v8_CY273Z  sky130_fd_pr__nfet_01v8_CY273Z_1
timestamp 1668290293
transform 0 1 58490 -1 0 147676
box -496 -260 496 260
use sky130_fd_pr__nfet_01v8_CY273Z  sky130_fd_pr__nfet_01v8_CY273Z_2
timestamp 1668290293
transform 0 1 59010 -1 0 147676
box -496 -260 496 260
use sky130_fd_pr__nfet_01v8_CY273Z  sky130_fd_pr__nfet_01v8_CY273Z_3
timestamp 1668290293
transform 0 1 59530 -1 0 147676
box -496 -260 496 260
use sky130_fd_pr__nfet_01v8_DPBXBZ  sky130_fd_pr__nfet_01v8_DPBXBZ_0
timestamp 1668293870
transform 1 0 554859 0 1 152234
box -783 -710 783 710
use sky130_fd_pr__nfet_01v8_SBZDCA  sky130_fd_pr__nfet_01v8_SBZDCA_0
timestamp 1669386980
transform 1 0 556317 0 1 152234
box -263 -710 263 710
use sky130_fd_pr__nfet_01v8_UBS3CQ  sky130_fd_pr__nfet_01v8_UBS3CQ_0
timestamp 1668293870
transform 0 1 553822 -1 0 151915
box -321 -260 321 260
use sky130_fd_pr__nfet_01v8_UBS3CQ  sky130_fd_pr__nfet_01v8_UBS3CQ_1
timestamp 1668293870
transform 0 1 553822 -1 0 152557
box -321 -260 321 260
use sky130_fd_pr__pfet_01v8_A7FR94  sky130_fd_pr__pfet_01v8_A7FR94_0
timestamp 1668293870
transform 0 1 553894 -1 0 153444
box -321 -319 321 319
use sky130_fd_pr__pfet_01v8_A7FR94  sky130_fd_pr__pfet_01v8_A7FR94_1
timestamp 1668293870
transform 0 1 553894 -1 0 154086
box -321 -319 321 319
use sky130_fd_pr__pfet_01v8_UJR9GH  sky130_fd_pr__pfet_01v8_UJR9GH_0
timestamp 1669386980
transform 1 0 556269 0 1 153825
box -455 -719 455 719
use sky130_fd_pr__pfet_01v8_YKSYY8  sky130_fd_pr__pfet_01v8_YKSYY8_0
timestamp 1668293870
transform 1 0 554839 0 1 153827
box -629 -719 629 719
use sky130_fd_pr__res_xhigh_po_5p73_2AHZHE  sky130_fd_pr__res_xhigh_po_5p73_2AHZHE_1
timestamp 1668288961
transform 0 1 58372 -1 0 128325
box -1981 -5102 1981 5102
use sky130_fd_pr__res_xhigh_po_5p73_2AHZHE  sky130_fd_pr__res_xhigh_po_5p73_2AHZHE_2
timestamp 1668288961
transform 0 1 58372 -1 0 124363
box -1981 -5102 1981 5102
use sky130_fd_pr__res_xhigh_po_5p73_2AHZHE  sky130_fd_pr__res_xhigh_po_5p73_2AHZHE_3
timestamp 1668288961
transform 0 1 58372 -1 0 120401
box -1981 -5102 1981 5102
use sky130_fd_pr__res_xhigh_po_5p73_2AHZHE  sky130_fd_pr__res_xhigh_po_5p73_2AHZHE_4
timestamp 1668288961
transform 0 1 58372 -1 0 116439
box -1981 -5102 1981 5102
use switched_cap  switched_cap_0
timestamp 1667842615
transform -1 0 358010 0 -1 391814
box -6253 -57972 42538 2189
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
