magic
tech sky130A
magscale 1 2
timestamp 1665942972
<< locali >>
rect -425 1474 -329 1508
rect 381 1474 897 1508
rect 1607 1474 1705 1508
rect -425 1412 -391 1474
rect -391 1032 -277 1330
rect -425 888 -391 950
rect 443 888 477 1474
rect 803 1330 837 1474
rect 803 1306 951 1330
rect 837 1052 951 1306
rect 803 1032 951 1052
rect 1671 1032 1705 1474
rect 803 888 837 1032
rect 1671 998 2643 1032
rect 3815 998 3977 1032
rect 1671 888 1705 998
rect -425 854 1705 888
rect -19 738 77 772
rect 625 738 893 772
rect 1441 738 1538 772
rect -19 678 15 738
rect -423 644 -327 678
rect -189 644 15 678
rect -423 582 -389 644
rect -423 -236 -389 122
rect -423 -740 -389 -678
rect -127 582 15 644
rect -93 116 15 582
rect -127 -118 15 116
rect 689 676 830 738
rect 723 -24 830 676
rect 1504 676 1538 738
rect 1504 150 1505 676
rect 1503 130 1505 150
rect 1539 130 1707 150
rect 1503 116 1707 130
rect 2257 116 2353 150
rect 689 -118 830 -24
rect 1504 -20 1645 116
rect 2319 54 2353 116
rect 1504 -118 1759 -20
rect -127 -260 1759 -118
rect -127 -740 15 -260
rect 689 -396 830 -260
rect 1504 -396 1759 -260
rect 575 -604 830 -396
rect 1389 -604 1759 -396
rect 689 -740 830 -604
rect 1504 -740 1645 -604
rect 2319 -740 2353 -678
rect -423 -774 -327 -740
rect -189 -774 77 -740
rect 597 -774 995 -740
rect 1353 -774 1765 -740
rect 2197 -774 2353 -740
rect 2435 -740 2469 998
rect 3943 -740 3977 998
rect 2435 -774 3977 -740
<< viali >>
rect -329 1474 381 1508
rect 897 1474 1607 1508
rect -425 950 -391 1412
rect 803 1052 837 1306
rect 2643 998 3815 1032
rect 77 738 625 772
rect 893 738 1441 772
rect -327 644 -189 678
rect -423 122 -389 582
rect -423 -678 -389 -236
rect -127 116 -93 582
rect 689 -24 723 676
rect 1505 130 1539 676
rect 1707 116 2257 150
rect 2319 -678 2353 54
rect -327 -774 -189 -740
rect 77 -774 597 -740
rect 995 -774 1353 -740
rect 1765 -774 2197 -740
<< metal1 >>
rect 1951 1682 2435 1692
rect 1951 1582 1961 1682
rect 2425 1582 2435 1682
rect -439 1462 -335 1520
rect 383 1462 897 1520
rect 1609 1462 1715 1520
rect -439 1412 -379 1462
rect -439 950 -425 1412
rect -391 1330 -379 1412
rect -265 1366 1545 1422
rect 1951 1408 2435 1582
rect -391 1314 -271 1330
rect -189 1320 -143 1366
rect 67 1320 113 1366
rect 323 1320 369 1366
rect -391 1048 -329 1314
rect -277 1048 -271 1314
rect -391 1032 -271 1048
rect -199 1314 -133 1320
rect -199 1048 -193 1314
rect -139 1048 -133 1314
rect -199 1042 -133 1048
rect -67 1314 -9 1320
rect -67 1048 -65 1314
rect -11 1048 -9 1314
rect -67 1042 -9 1048
rect 57 1314 123 1320
rect 57 1048 63 1314
rect 117 1048 123 1314
rect 57 1042 123 1048
rect 189 1314 247 1320
rect 189 1048 191 1314
rect 245 1048 247 1314
rect 189 1042 247 1048
rect 313 1314 379 1320
rect 313 1048 319 1314
rect 373 1048 379 1314
rect 313 1042 379 1048
rect 779 1314 957 1330
rect 779 1306 899 1314
rect 779 1052 803 1306
rect 837 1052 899 1306
rect 779 1048 899 1052
rect 951 1048 957 1314
rect -391 950 -379 1032
rect -189 996 -143 1042
rect 67 996 113 1042
rect 323 998 369 1042
rect 779 1032 957 1048
rect 1029 1314 1095 1320
rect 1029 1048 1035 1314
rect 1089 1048 1095 1314
rect 1029 1042 1095 1048
rect 1157 1314 1223 1320
rect 1157 1048 1163 1314
rect 1217 1048 1223 1314
rect 1157 1042 1223 1048
rect 1285 1314 1351 1320
rect 1285 1048 1291 1314
rect 1345 1048 1351 1314
rect 1285 1042 1351 1048
rect 1413 1314 1479 1320
rect 1413 1048 1419 1314
rect 1473 1048 1479 1314
rect 1413 1042 1479 1048
rect 1541 1314 1607 1320
rect 1541 1048 1547 1314
rect 1601 1048 1607 1314
rect 1541 1042 1607 1048
rect 1859 1204 2435 1408
rect 304 996 369 998
rect -439 840 -379 950
rect -265 940 1545 996
rect 1859 946 2343 1204
rect 2631 1042 3831 1044
rect 2631 988 2643 1042
rect 3815 988 3831 1042
rect 1767 890 3816 946
rect 1767 876 1823 890
rect 1767 814 1823 820
rect -135 772 1545 780
rect -135 738 77 772
rect 625 738 893 772
rect 1441 738 1545 772
rect -135 730 1545 738
rect -135 684 -85 730
rect -429 678 -85 684
rect -429 644 -327 678
rect -189 644 -85 678
rect -429 638 -85 644
rect -429 582 -381 638
rect -429 122 -423 582
rect -389 122 -381 582
rect -135 582 -85 638
rect -291 532 -227 538
rect -291 132 -285 532
rect -233 132 -227 532
rect -291 126 -227 132
rect -429 110 -381 122
rect -135 116 -127 582
rect -93 116 -85 582
rect -135 104 -85 116
rect 3 630 481 686
rect 677 676 735 730
rect 3 40 53 630
rect -459 -10 53 40
rect 81 586 149 592
rect 81 34 87 586
rect 143 34 149 586
rect 81 28 149 34
rect 177 586 241 592
rect 177 34 183 586
rect 235 34 241 586
rect 177 28 241 34
rect 271 586 339 592
rect 271 34 277 586
rect 333 34 339 586
rect 271 28 339 34
rect 367 586 431 592
rect 367 34 373 586
rect 425 34 431 586
rect 367 28 431 34
rect 463 586 531 592
rect 463 34 469 586
rect 525 34 531 586
rect 463 28 531 34
rect 563 586 627 592
rect 563 34 569 586
rect 621 34 627 586
rect 563 28 627 34
rect -459 -50 577 -10
rect 677 -24 689 676
rect 723 -24 735 676
rect 677 -36 735 -24
rect 807 630 1295 686
rect 1497 676 1545 730
rect 807 -10 863 630
rect 893 586 957 592
rect 893 34 899 586
rect 951 34 957 586
rect 893 22 957 34
rect 989 586 1053 592
rect 989 34 995 586
rect 1047 34 1053 586
rect 989 28 1053 34
rect 1083 586 1147 592
rect 1083 34 1089 586
rect 1141 34 1147 586
rect 1083 22 1147 34
rect 1183 586 1247 592
rect 1183 34 1189 586
rect 1241 34 1247 586
rect 1183 28 1247 34
rect 1279 586 1343 592
rect 1279 34 1285 586
rect 1337 34 1343 586
rect 1279 22 1343 34
rect 1375 586 1439 592
rect 1375 34 1381 586
rect 1433 34 1439 586
rect 1497 130 1505 676
rect 1539 156 1545 676
rect 1539 150 2363 156
rect 1539 130 1707 150
rect 1497 116 1707 130
rect 2257 116 2363 150
rect 1497 106 2363 116
rect 1375 28 1439 34
rect 1549 8 2111 64
rect 2311 54 2363 106
rect 3 -66 577 -50
rect 807 -66 1391 -10
rect 807 -94 899 -66
rect -459 -186 899 -94
rect -437 -236 -373 -224
rect -437 -678 -423 -236
rect -389 -678 -373 -236
rect 1549 -312 1605 8
rect 83 -368 1605 -312
rect 83 -400 135 -368
rect -293 -600 135 -400
rect 175 -412 241 -406
rect 175 -588 181 -412
rect 235 -588 241 -412
rect 175 -594 241 -588
rect -437 -724 -373 -678
rect 83 -632 135 -600
rect 281 -632 327 -368
rect 367 -412 433 -406
rect 367 -588 373 -412
rect 427 -588 433 -412
rect 367 -594 433 -588
rect 473 -632 519 -368
rect 559 -412 625 -406
rect 559 -588 565 -412
rect 619 -588 625 -412
rect 559 -594 625 -588
rect 735 -632 783 -368
rect 893 -412 957 -406
rect 893 -588 899 -412
rect 951 -588 957 -412
rect 893 -594 957 -588
rect 989 -412 1055 -406
rect 989 -588 995 -412
rect 1049 -588 1055 -412
rect 989 -594 1055 -588
rect 1087 -412 1151 -406
rect 1087 -588 1093 -412
rect 1145 -588 1151 -412
rect 1087 -594 1151 -588
rect 1183 -412 1249 -406
rect 1183 -588 1189 -412
rect 1241 -588 1249 -412
rect 1183 -594 1249 -588
rect 1279 -412 1343 -406
rect 1279 -588 1285 -412
rect 1337 -588 1343 -412
rect 1279 -594 1343 -588
rect 1375 -412 1439 -406
rect 1375 -588 1381 -412
rect 1433 -588 1439 -412
rect 1375 -594 1439 -588
rect 1549 -632 1605 -368
rect 1707 -36 1771 -30
rect 1707 -588 1713 -36
rect 1765 -588 1771 -36
rect 1707 -594 1771 -588
rect 1807 -36 1871 -30
rect 1807 -588 1813 -36
rect 1865 -588 1871 -36
rect 1807 -594 1871 -588
rect 1903 -36 1967 -30
rect 1903 -588 1909 -36
rect 1961 -588 1967 -36
rect 1903 -594 1967 -588
rect 1999 -36 2063 -30
rect 1999 -588 2005 -36
rect 2057 -588 2063 -36
rect 1999 -594 2063 -588
rect 2095 -36 2159 -30
rect 2095 -588 2101 -36
rect 2153 -588 2159 -36
rect 2095 -594 2159 -588
rect 2191 -36 2255 -30
rect 2191 -588 2197 -36
rect 2249 -588 2255 -36
rect 2191 -594 2255 -588
rect 83 -688 2207 -632
rect 2311 -678 2319 54
rect 2353 -678 2363 54
rect -437 -730 605 -724
rect -437 -740 241 -730
rect -437 -774 -327 -740
rect -189 -774 77 -740
rect -437 -782 241 -774
rect 597 -782 605 -730
rect -437 -788 605 -782
rect 989 -730 1359 -724
rect 2311 -726 2363 -678
rect 2397 -632 2453 890
rect 2531 838 2595 844
rect 2531 -580 2537 838
rect 2589 -580 2595 838
rect 2531 -586 2595 -580
rect 2661 838 2725 844
rect 2661 -580 2667 838
rect 2719 -580 2725 838
rect 2661 -586 2725 -580
rect 2791 838 2855 844
rect 2791 -580 2797 838
rect 2849 -580 2855 838
rect 2791 -586 2855 -580
rect 2917 838 2981 844
rect 2917 -580 2923 838
rect 2975 -580 2981 838
rect 2917 -586 2981 -580
rect 3047 838 3111 844
rect 3047 -580 3053 838
rect 3105 -580 3111 838
rect 3047 -586 3111 -580
rect 3173 838 3237 844
rect 3173 -580 3179 838
rect 3231 -580 3237 838
rect 3173 -586 3237 -580
rect 3303 838 3367 844
rect 3303 -580 3309 838
rect 3361 -580 3367 838
rect 3303 -586 3367 -580
rect 3429 838 3493 844
rect 3429 -580 3435 838
rect 3487 -580 3493 838
rect 3429 -586 3493 -580
rect 3559 838 3623 844
rect 3559 -580 3565 838
rect 3617 -580 3623 838
rect 3559 -586 3623 -580
rect 3685 838 3749 844
rect 3685 -580 3691 838
rect 3743 -580 3749 838
rect 3685 -586 3749 -580
rect 3815 838 3879 844
rect 3815 -580 3821 838
rect 3873 -580 3879 838
rect 3815 -586 3879 -580
rect 2397 -688 3816 -632
rect 989 -782 995 -730
rect 1353 -782 1359 -730
rect 989 -788 1359 -782
rect 1759 -732 2363 -726
rect 1759 -786 1765 -732
rect 2197 -786 2363 -732
rect 1759 -792 2363 -786
<< via1 >>
rect 1961 1582 2425 1682
rect -335 1508 383 1520
rect -335 1474 -329 1508
rect -329 1474 381 1508
rect 381 1474 383 1508
rect -335 1462 383 1474
rect 897 1508 1609 1520
rect 897 1474 1607 1508
rect 1607 1474 1609 1508
rect 897 1462 1609 1474
rect -329 1048 -277 1314
rect -193 1048 -139 1314
rect -65 1048 -11 1314
rect 63 1048 117 1314
rect 191 1048 245 1314
rect 319 1048 373 1314
rect 899 1048 951 1314
rect 1035 1048 1089 1314
rect 1163 1048 1217 1314
rect 1291 1048 1345 1314
rect 1419 1048 1473 1314
rect 1547 1048 1601 1314
rect 2643 1032 3815 1042
rect 2643 998 3815 1032
rect 2643 988 3815 998
rect 1767 820 1823 876
rect -285 132 -233 532
rect 87 34 143 586
rect 183 34 235 586
rect 277 34 333 586
rect 373 34 425 586
rect 469 34 525 586
rect 569 34 621 586
rect 899 34 951 586
rect 995 34 1047 586
rect 1089 34 1141 586
rect 1189 34 1241 586
rect 1285 34 1337 586
rect 1381 34 1433 586
rect 181 -588 235 -412
rect 373 -588 427 -412
rect 565 -588 619 -412
rect 899 -588 951 -412
rect 995 -588 1049 -412
rect 1093 -588 1145 -412
rect 1189 -588 1241 -412
rect 1285 -588 1337 -412
rect 1381 -588 1433 -412
rect 1713 -588 1765 -36
rect 1813 -588 1865 -36
rect 1909 -588 1961 -36
rect 2005 -588 2057 -36
rect 2101 -588 2153 -36
rect 2197 -588 2249 -36
rect 241 -740 597 -730
rect 241 -774 597 -740
rect 241 -782 597 -774
rect 2537 -580 2589 838
rect 2667 -580 2719 838
rect 2797 -580 2849 838
rect 2923 -580 2975 838
rect 3053 -580 3105 838
rect 3179 -580 3231 838
rect 3309 -580 3361 838
rect 3435 -580 3487 838
rect 3565 -580 3617 838
rect 3691 -580 3743 838
rect 3821 -580 3873 838
rect 995 -740 1353 -730
rect 995 -774 1353 -740
rect 995 -782 1353 -774
rect 1765 -740 2197 -732
rect 1765 -774 2197 -740
rect 1765 -786 2197 -774
<< metal2 >>
rect 1951 1682 2435 1692
rect 1951 1582 1961 1682
rect 2425 1582 2435 1682
rect 1951 1574 2435 1582
rect -335 1520 1741 1544
rect 383 1462 897 1520
rect 1609 1462 1741 1520
rect -335 1452 1741 1462
rect -335 1314 -271 1452
rect -335 1048 -329 1314
rect -277 1048 -271 1314
rect -335 738 -271 1048
rect -199 1314 -133 1320
rect -199 1048 -193 1314
rect -139 1048 -133 1314
rect -199 910 -133 1048
rect -67 1314 -9 1452
rect -67 1048 -65 1314
rect -11 1048 -9 1314
rect -67 1042 -9 1048
rect 57 1314 123 1320
rect 57 1048 63 1314
rect 117 1048 123 1314
rect 57 910 123 1048
rect 189 1314 247 1452
rect 189 1048 191 1314
rect 245 1048 247 1314
rect 189 1042 247 1048
rect 313 1314 379 1320
rect 313 1048 319 1314
rect 373 1048 379 1314
rect 313 910 379 1048
rect 893 1314 957 1452
rect 893 1048 899 1314
rect 951 1048 957 1314
rect 893 1042 957 1048
rect 1029 1314 1095 1320
rect 1029 1048 1035 1314
rect 1089 1048 1095 1314
rect 1029 910 1095 1048
rect 1161 1314 1219 1452
rect 1161 1048 1163 1314
rect 1217 1048 1219 1314
rect 1161 1042 1219 1048
rect 1285 1314 1351 1320
rect 1285 1048 1291 1314
rect 1345 1048 1351 1314
rect 1285 910 1351 1048
rect 1417 1314 1475 1452
rect 1417 1048 1419 1314
rect 1473 1048 1475 1314
rect 1417 1042 1475 1048
rect 1541 1314 1607 1320
rect 1541 1048 1547 1314
rect 1601 1048 1607 1314
rect 1541 910 1607 1048
rect 1649 1144 1741 1452
rect 3007 1144 3607 1614
rect 1649 1042 4013 1144
rect 1649 988 2643 1042
rect 3815 988 4013 1042
rect 1649 970 4013 988
rect -199 818 531 910
rect 1029 888 1607 910
rect -335 674 -227 738
rect -291 532 -227 674
rect -291 132 -285 532
rect -233 132 -227 532
rect -291 126 -227 132
rect 81 586 149 818
rect 81 34 87 586
rect 143 34 149 586
rect 81 28 149 34
rect 177 586 241 592
rect 177 34 183 586
rect 235 34 241 586
rect 177 -70 241 34
rect 271 586 339 818
rect 271 34 277 586
rect 333 34 339 586
rect 271 28 339 34
rect 367 586 431 592
rect 367 34 373 586
rect 425 34 431 586
rect 367 -70 431 34
rect 463 586 531 818
rect 989 878 1607 888
rect 989 876 1829 878
rect 989 820 1767 876
rect 1823 820 1829 876
rect 989 818 1829 820
rect 2531 838 2595 844
rect 463 34 469 586
rect 525 34 531 586
rect 463 28 531 34
rect 563 586 627 592
rect 563 34 569 586
rect 621 34 627 586
rect 563 -70 627 34
rect 893 586 957 592
rect 893 34 899 586
rect 951 34 957 586
rect 893 -70 957 34
rect 989 586 1053 818
rect 989 34 995 586
rect 1047 34 1053 586
rect 989 28 1053 34
rect 1083 586 1147 592
rect 1083 34 1089 586
rect 1141 34 1147 586
rect 1083 -70 1147 34
rect 1183 586 1247 818
rect 1183 34 1189 586
rect 1241 34 1247 586
rect 1183 28 1247 34
rect 1279 586 1343 592
rect 1279 34 1285 586
rect 1337 34 1343 586
rect 1279 -70 1343 34
rect 1375 586 1439 818
rect 1375 34 1381 586
rect 1433 34 1439 586
rect 1375 28 1439 34
rect 1807 62 2471 186
rect 177 -134 1343 -70
rect 175 -412 241 -406
rect 175 -588 181 -412
rect 235 -588 241 -412
rect 175 -720 241 -588
rect 367 -412 433 -406
rect 367 -588 373 -412
rect 427 -588 433 -412
rect 367 -720 433 -588
rect 559 -412 625 -406
rect 559 -588 565 -412
rect 619 -588 625 -412
rect 559 -720 625 -588
rect 893 -412 957 -134
rect 893 -588 899 -412
rect 951 -588 957 -412
rect 893 -594 957 -588
rect 989 -412 1055 -406
rect 989 -588 995 -412
rect 1049 -588 1055 -412
rect 989 -720 1055 -588
rect 1087 -412 1151 -134
rect 1087 -588 1093 -412
rect 1145 -588 1151 -412
rect 1087 -594 1151 -588
rect 1183 -412 1249 -406
rect 1183 -588 1189 -412
rect 1241 -588 1249 -412
rect 1183 -720 1249 -588
rect 1279 -412 1343 -134
rect 1707 -36 1771 -30
rect 1279 -588 1285 -412
rect 1337 -588 1343 -412
rect 1279 -594 1343 -588
rect 1375 -412 1439 -406
rect 1375 -588 1381 -412
rect 1433 -588 1439 -412
rect 1375 -720 1439 -588
rect 1707 -588 1713 -36
rect 1765 -588 1771 -36
rect 1707 -720 1771 -588
rect 1807 -36 1871 62
rect 1807 -588 1813 -36
rect 1865 -588 1871 -36
rect 1807 -594 1871 -588
rect 1903 -36 1967 -30
rect 1903 -588 1909 -36
rect 1961 -588 1967 -36
rect 1903 -720 1967 -588
rect 1999 -36 2063 62
rect 1999 -588 2005 -36
rect 2057 -588 2063 -36
rect 1999 -594 2063 -588
rect 2095 -36 2159 -30
rect 2095 -588 2101 -36
rect 2153 -588 2159 -36
rect 2095 -720 2159 -588
rect 2191 -36 2255 62
rect 2191 -588 2197 -36
rect 2249 -588 2255 -36
rect 2191 -594 2255 -588
rect 2347 -688 2471 62
rect 2531 -580 2537 838
rect 2589 -580 2595 838
rect 2531 -688 2595 -580
rect 2661 838 2725 970
rect 2661 -580 2667 838
rect 2719 -580 2725 838
rect 2661 -586 2725 -580
rect 2791 838 2855 844
rect 2791 -580 2797 838
rect 2849 -580 2855 838
rect 2791 -688 2855 -580
rect 2917 838 2981 970
rect 2917 -580 2923 838
rect 2975 -580 2981 838
rect 2917 -586 2981 -580
rect 3047 838 3111 844
rect 3047 -580 3053 838
rect 3105 -580 3111 838
rect 3047 -688 3111 -580
rect 3173 838 3237 970
rect 3173 -580 3179 838
rect 3231 -580 3237 838
rect 3173 -586 3237 -580
rect 3303 838 3367 844
rect 3303 -580 3309 838
rect 3361 -580 3367 838
rect 3303 -688 3367 -580
rect 3429 838 3493 970
rect 3429 -580 3435 838
rect 3487 -580 3493 838
rect 3429 -586 3493 -580
rect 3559 838 3623 844
rect 3559 -580 3565 838
rect 3617 -580 3623 838
rect 3559 -688 3623 -580
rect 3685 838 3749 970
rect 3685 -580 3691 838
rect 3743 -580 3749 838
rect 3685 -586 3749 -580
rect 3815 838 3879 844
rect 3815 -580 3821 838
rect 3873 -580 3879 838
rect 3815 -688 3879 -580
rect 175 -730 2237 -720
rect 175 -782 241 -730
rect 597 -782 995 -730
rect 1353 -732 2237 -730
rect 1353 -782 1765 -732
rect 175 -786 1765 -782
rect 2197 -786 2237 -732
rect 175 -810 2237 -786
rect 2347 -792 3879 -688
rect 1619 -952 2219 -810
rect 2347 -812 2571 -792
rect 2561 -944 2571 -812
rect 3673 -812 3879 -792
rect 3673 -944 3681 -812
rect 2561 -954 3681 -944
<< via2 >>
rect 1961 1582 2425 1682
rect 2571 -944 3673 -792
<< metal3 >>
rect 1951 1682 2435 1692
rect 1951 1582 1961 1682
rect 2425 1582 2435 1682
rect 1951 1386 2435 1582
rect 2561 -792 3681 -784
rect 2561 -944 2571 -792
rect 3673 -944 3681 -792
rect 2561 -954 3681 -944
<< via3 >>
rect 1961 1582 2425 1682
rect 2571 -944 3673 -792
<< metal4 >>
rect 1951 1996 2711 2020
rect 1951 1724 1975 1996
rect 2687 1724 2711 1996
rect 1951 1682 2711 1724
rect 1951 1582 1961 1682
rect 2425 1582 2711 1682
rect 1951 1576 2711 1582
rect 2561 -792 3681 -684
rect 2561 -944 2571 -792
rect 3673 -944 3681 -792
rect 2561 -954 3681 -944
<< via4 >>
rect 1975 1724 2687 1996
<< metal5 >>
rect 1951 1996 2711 2020
rect 1951 1724 1975 1996
rect 2687 1724 2711 1996
rect 1951 1378 2711 1724
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_0
timestamp 1665661446
transform -1 0 2656 0 -1 396
box -1150 -1100 1049 1100
use sky130_fd_pr__cap_mim_m3_2_6ZNTNB  sky130_fd_pr__cap_mim_m3_2_6ZNTNB_0
timestamp 1665661005
transform 1 0 2959 0 1 394
box -1351 -1100 849 1100
use sky130_fd_pr__nfet_01v8_lvt_46VND8  sky130_fd_pr__nfet_01v8_lvt_46VND8_0
timestamp 1665942972
transform 1 0 1982 0 1 -312
box -407 -498 407 498
use sky130_fd_pr__nfet_01v8_lvt_46VND8  sky130_fd_pr__nfet_01v8_lvt_46VND8_1
timestamp 1665942972
transform 1 0 352 0 1 310
box -407 -498 407 498
use sky130_fd_pr__nfet_01v8_lvt_46VND8  sky130_fd_pr__nfet_01v8_lvt_46VND8_2
timestamp 1665942972
transform 1 0 1167 0 1 310
box -407 -498 407 498
use sky130_fd_pr__nfet_01v8_lvt_595QY5  sky130_fd_pr__nfet_01v8_lvt_595QY5_0
timestamp 1665942907
transform 1 0 352 0 1 -500
box -407 -310 407 310
use sky130_fd_pr__nfet_01v8_lvt_595QY5  sky130_fd_pr__nfet_01v8_lvt_595QY5_1
timestamp 1665942907
transform 1 0 1167 0 1 -500
box -407 -310 407 310
use sky130_fd_pr__pfet_01v8_lvt_4YVKJ3  sky130_fd_pr__pfet_01v8_lvt_4YVKJ3_0
timestamp 1665942722
transform 1 0 26 0 1 1181
box -487 -363 487 363
use sky130_fd_pr__pfet_01v8_lvt_4YVKJ3  sky130_fd_pr__pfet_01v8_lvt_4YVKJ3_1
timestamp 1665942722
transform 1 0 1254 0 1 1181
box -487 -363 487 363
use sky130_fd_pr__pfet_01v8_lvt_MUFCUN  sky130_fd_pr__pfet_01v8_lvt_MUFCUN_1
timestamp 1665678605
transform 1 0 3207 0 1 129
box -807 -939 807 939
use sky130_fd_pr__res_xhigh_po_0p35_NZJDJZ  sky130_fd_pr__res_xhigh_po_0p35_NZJDJZ_0
timestamp 1665674792
transform 1 0 -258 0 1 -48
box -201 -762 201 762
<< labels >>
rlabel metal1 -447 -14 -447 -14 3 Inv
port 1 e
rlabel metal2 1929 -928 1931 -928 5 Vss
port 5 s
rlabel metal2 3279 1588 3279 1588 1 Vdd
port 4 n
rlabel metal4 2845 -948 2845 -948 5 Out
port 3 s
rlabel metal1 -445 -140 -445 -140 7 NonInv
port 2 w
<< end >>
