magic
tech sky130A
magscale 1 2
timestamp 1668785164
<< obsactive >>
rect -74 5994 6226 7172
rect -74 304 818 5994
rect 5334 304 6226 5994
rect -74 -306 6226 304
rect -74 -5996 818 -306
rect 5334 -5996 6226 -306
rect -74 -6606 6226 -5996
rect -74 -12296 818 -6606
rect 5334 -12296 6226 -6606
rect -74 -12906 6226 -12296
rect -74 -18596 818 -12906
rect 5334 -18596 6226 -12906
rect -74 -19206 6226 -18596
rect -74 -24896 818 -19206
rect 5334 -24896 6226 -19206
rect -74 -25506 6226 -24896
rect -74 -31196 818 -25506
rect 5334 -31196 6226 -25506
rect -74 -31806 6226 -31196
rect -74 -37496 818 -31806
rect 5334 -37496 6226 -31806
rect -74 -38106 6226 -37496
rect -74 -43796 818 -38106
rect 5334 -43796 6226 -38106
rect -74 -44406 6226 -43796
rect -74 -50096 818 -44406
rect 5334 -50096 6226 -44406
rect -74 -50706 6226 -50096
rect -74 -56396 818 -50706
rect 5334 -56396 6226 -50706
rect -74 -57006 6226 -56396
rect -74 -62696 818 -57006
rect 5334 -62696 6226 -57006
rect -74 -63306 6226 -62696
rect -74 -68996 818 -63306
rect 5334 -68996 6226 -63306
rect -74 -69606 6226 -68996
rect -74 -75296 818 -69606
rect 5334 -75296 6226 -69606
rect -74 -75906 6226 -75296
rect -74 -81596 818 -75906
rect 5334 -81596 6226 -75906
rect -74 -82206 6226 -81596
rect -74 -87896 818 -82206
rect 5334 -87896 6226 -82206
rect -74 -88506 6226 -87896
rect -74 -94196 818 -88506
rect 5334 -94196 6226 -88506
rect -74 -94806 6226 -94196
rect -74 -100496 818 -94806
rect 5334 -100496 6226 -94806
rect -74 -101106 6226 -100496
rect -74 -106796 818 -101106
rect 5334 -106796 6226 -101106
rect -74 -107406 6226 -106796
rect -74 -113096 818 -107406
rect 5334 -113096 6226 -107406
rect -74 -113706 6226 -113096
rect -74 -119396 818 -113706
rect 5334 -119396 6226 -113706
rect -74 -120006 6226 -119396
rect -74 -125696 818 -120006
rect 5334 -125696 6226 -120006
rect -74 -126306 6226 -125696
rect -74 -131996 818 -126306
rect 5334 -131996 6226 -126306
rect -74 -132606 6226 -131996
rect -74 -138296 818 -132606
rect 5334 -138296 6226 -132606
rect -74 -138906 6226 -138296
rect -74 -144596 818 -138906
rect 5334 -144596 6226 -138906
rect -74 -145206 6226 -144596
rect -74 -150896 818 -145206
rect 5334 -150896 6226 -145206
rect -74 -151506 6226 -150896
rect -74 -157196 818 -151506
rect 5334 -157196 6226 -151506
rect -74 -157806 6226 -157196
rect -74 -163496 818 -157806
rect 5334 -163496 6226 -157806
rect -74 -164106 6226 -163496
rect -74 -169796 818 -164106
rect 5334 -169796 6226 -164106
rect -74 -170406 6226 -169796
rect -74 -176096 818 -170406
rect 5334 -176096 6226 -170406
rect -74 -176706 6226 -176096
rect -74 -182396 818 -176706
rect 5334 -182396 6226 -176706
rect -74 -183006 6226 -182396
rect -74 -188696 818 -183006
rect 5334 -188696 6226 -183006
rect -74 -189306 6226 -188696
rect -74 -194996 818 -189306
rect 5334 -194996 6226 -189306
rect -74 -196225 6226 -194996
<< metal1 >>
rect 1176 6854 1576 6874
rect 1176 6594 1196 6854
rect 1556 6594 1576 6854
rect 1176 6274 1576 6594
rect 4575 6854 4975 6874
rect 4575 6594 4595 6854
rect 4955 6594 4975 6854
rect 4575 6274 4975 6594
rect 1176 6074 4975 6274
rect 1176 -195126 1376 6074
rect 4775 -195126 4975 6074
rect 1176 -195326 4975 -195126
rect 1176 -195646 1577 -195326
rect 1176 -195906 1197 -195646
rect 1557 -195906 1577 -195646
rect 1176 -195926 1577 -195906
rect 4576 -195646 4975 -195326
rect 4576 -195906 4596 -195646
rect 4955 -195906 4975 -195646
rect 4576 -195926 4975 -195906
<< via1 >>
rect 1196 6594 1556 6854
rect 4595 6594 4955 6854
rect 1197 -195906 1557 -195646
rect 4596 -195906 4955 -195646
<< metal2 >>
rect 2776 7133 3376 7153
rect 1176 6854 1576 6874
rect 1176 6594 1196 6854
rect 1556 6594 1576 6854
rect 1176 6574 1576 6594
rect 2776 6773 2796 7133
rect 3356 6773 3376 7133
rect 2776 6424 3376 6773
rect 4575 6854 4975 6874
rect 4575 6594 4595 6854
rect 4955 6594 4975 6854
rect 4575 6574 4975 6594
rect 894 6274 5258 6424
rect 894 -195326 1044 6274
rect 5108 -195326 5258 6274
rect 894 -195476 5258 -195326
rect 1176 -195646 1577 -195626
rect 1176 -195906 1197 -195646
rect 1557 -195906 1577 -195646
rect 1176 -195926 1577 -195906
rect 2776 -195825 3376 -195476
rect 2776 -196185 2796 -195825
rect 3356 -196185 3376 -195825
rect 4576 -195646 4975 -195626
rect 4576 -195906 4596 -195646
rect 4955 -195906 4975 -195646
rect 4576 -195926 4975 -195906
rect 2776 -196205 3376 -196185
<< via2 >>
rect 1196 6594 1556 6854
rect 2796 6773 3356 7133
rect 4595 6594 4955 6854
rect 1197 -195906 1557 -195646
rect 2796 -196185 3356 -195825
rect 4596 -195906 4955 -195646
<< metal3 >>
rect 2751 7133 3394 7173
rect 1176 6854 1576 6874
rect 1176 6594 1196 6854
rect 1556 6594 1576 6854
rect 1176 6574 1576 6594
rect 2751 6773 2796 7133
rect 3356 6773 3394 7133
rect 2751 6084 3394 6773
rect 4575 6854 4975 6874
rect 4575 6594 4595 6854
rect 4955 6594 4975 6854
rect 4575 6574 4975 6594
rect 1176 -195646 1577 -195626
rect 1176 -195906 1197 -195646
rect 1557 -195906 1577 -195646
rect 1176 -195926 1577 -195906
rect 2758 -195825 3401 -195136
rect 2758 -196185 2796 -195825
rect 3356 -196185 3401 -195825
rect 4576 -195646 4975 -195626
rect 4576 -195906 4596 -195646
rect 4955 -195906 4975 -195646
rect 4576 -195926 4975 -195906
rect 2758 -196225 3401 -196185
<< via3 >>
rect 1196 6594 1556 6854
rect 2796 6773 3356 7133
rect 4595 6594 4955 6854
rect 1197 -195906 1557 -195646
rect 2796 -196185 3356 -195825
rect 4596 -195906 4955 -195646
<< metal4 >>
rect 2776 7133 3376 7153
rect 1176 6854 1576 6874
rect 1176 6594 1196 6854
rect 1556 6594 1576 6854
rect 2776 6773 2796 7133
rect 3356 6773 3376 7133
rect 2776 6753 3376 6773
rect 4575 6854 4975 6874
rect 1176 6108 1576 6594
rect 4575 6594 4595 6854
rect 4955 6594 4975 6854
rect 4575 6108 4975 6594
rect 1176 -195646 1577 -195160
rect 1176 -195906 1197 -195646
rect 1557 -195906 1577 -195646
rect 4576 -195646 4975 -195160
rect 1176 -195926 1577 -195906
rect 2776 -195825 3376 -195805
rect 2776 -196185 2796 -195825
rect 3356 -196185 3376 -195825
rect 4576 -195906 4596 -195646
rect 4955 -195906 4975 -195646
rect 4576 -195926 4975 -195906
rect 2776 -196205 3376 -196185
<< via4 >>
rect 2796 6773 3356 7133
rect 2796 -196185 3356 -195825
<< metal5 >>
rect 2751 7133 3394 7173
rect 2751 6773 2796 7133
rect 3356 6773 3394 7133
rect 2751 6084 3394 6773
rect 2758 -195825 3401 -195136
rect 2758 -196185 2796 -195825
rect 3356 -196185 3401 -195825
rect 2758 -196225 3401 -196185
use sky130_fd_pr__cap_mim_m3_1_U59KTN  sky130_fd_pr__cap_mim_m3_1_U59KTN_0
timestamp 1667066906
transform 1 0 3126 0 1 -94526
box -3200 -100800 3100 100800
use sky130_fd_pr__cap_mim_m3_2_U59KTN  sky130_fd_pr__cap_mim_m3_2_U59KTN_0
timestamp 1667067748
transform 1 0 3327 0 1 -94526
box -3401 -100800 2899 100800
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_0
timestamp 1667069478
transform 0 1 3076 -1 0 3149
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_1
timestamp 1667069478
transform 0 1 3076 -1 0 -3151
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_2
timestamp 1667069478
transform 0 1 3076 -1 0 -9451
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_3
timestamp 1667069478
transform 0 1 3076 -1 0 -15751
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_4
timestamp 1667069478
transform 0 1 3076 -1 0 -22051
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_5
timestamp 1667069478
transform 0 1 3076 -1 0 -28351
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_6
timestamp 1667069478
transform 0 1 3076 -1 0 -34651
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_7
timestamp 1667069478
transform 0 1 3076 -1 0 -40951
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_8
timestamp 1667069478
transform 0 1 3076 -1 0 -47251
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_9
timestamp 1667069478
transform 0 1 3076 -1 0 -53551
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_10
timestamp 1667069478
transform 0 1 3076 -1 0 -59851
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_11
timestamp 1667069478
transform 0 1 3076 -1 0 -66151
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_12
timestamp 1667069478
transform 0 1 3076 -1 0 -72451
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_13
timestamp 1667069478
transform 0 1 3076 -1 0 -78751
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_14
timestamp 1667069478
transform 0 1 3076 -1 0 -85051
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_15
timestamp 1667069478
transform 0 1 3076 -1 0 -91351
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_16
timestamp 1667069478
transform 0 1 3076 -1 0 -97651
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_17
timestamp 1667069478
transform 0 1 3076 -1 0 -103951
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_18
timestamp 1667069478
transform 0 1 3076 -1 0 -110251
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_19
timestamp 1667069478
transform 0 1 3076 -1 0 -116551
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_20
timestamp 1667069478
transform 0 1 3076 -1 0 -122851
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_21
timestamp 1667069478
transform 0 1 3076 -1 0 -129151
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_22
timestamp 1667069478
transform 0 1 3076 -1 0 -135451
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_23
timestamp 1667069478
transform 0 1 3076 -1 0 -141751
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_24
timestamp 1667069478
transform 0 1 3076 -1 0 -148051
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_25
timestamp 1667069478
transform 0 1 3076 -1 0 -154351
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_26
timestamp 1667069478
transform 0 1 3076 -1 0 -160651
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_27
timestamp 1667069478
transform 0 1 3076 -1 0 -166951
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_28
timestamp 1667069478
transform 0 1 3076 -1 0 -173251
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_29
timestamp 1667069478
transform 0 1 3076 -1 0 -179551
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_30
timestamp 1667069478
transform 0 1 3076 -1 0 -185851
box -2844 -2258 2844 2258
use sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ  sky130_fd_pr__nfet_g5v0d10v5_RTWZFQ_31
timestamp 1667069478
transform 0 1 3076 -1 0 -192151
box -2844 -2258 2844 2258
<< end >>
