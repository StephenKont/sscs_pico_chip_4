magic
tech sky130A
magscale 1 2
timestamp 1668293870
<< nwell >>
rect -629 -719 629 719
<< pmos >>
rect -433 -500 -183 500
rect -125 -500 125 500
rect 183 -500 433 500
<< pdiff >>
rect -491 488 -433 500
rect -491 -488 -479 488
rect -445 -488 -433 488
rect -491 -500 -433 -488
rect -183 488 -125 500
rect -183 -488 -171 488
rect -137 -488 -125 488
rect -183 -500 -125 -488
rect 125 488 183 500
rect 125 -488 137 488
rect 171 -488 183 488
rect 125 -500 183 -488
rect 433 488 491 500
rect 433 -488 445 488
rect 479 -488 491 488
rect 433 -500 491 -488
<< pdiffc >>
rect -479 -488 -445 488
rect -171 -488 -137 488
rect 137 -488 171 488
rect 445 -488 479 488
<< nsubdiff >>
rect -593 649 -497 683
rect 497 649 593 683
rect -593 587 -559 649
rect 559 587 593 649
rect -593 -649 -559 -587
rect 559 -649 593 -587
rect -593 -683 -497 -649
rect 497 -683 593 -649
<< nsubdiffcont >>
rect -497 649 497 683
rect -593 -587 -559 587
rect 559 -587 593 587
rect -497 -683 497 -649
<< poly >>
rect -433 581 -183 597
rect -433 547 -417 581
rect -199 547 -183 581
rect -433 500 -183 547
rect -125 581 125 597
rect -125 547 -109 581
rect 109 547 125 581
rect -125 500 125 547
rect 183 581 433 597
rect 183 547 199 581
rect 417 547 433 581
rect 183 500 433 547
rect -433 -547 -183 -500
rect -433 -581 -417 -547
rect -199 -581 -183 -547
rect -433 -597 -183 -581
rect -125 -547 125 -500
rect -125 -581 -109 -547
rect 109 -581 125 -547
rect -125 -597 125 -581
rect 183 -547 433 -500
rect 183 -581 199 -547
rect 417 -581 433 -547
rect 183 -597 433 -581
<< polycont >>
rect -417 547 -199 581
rect -109 547 109 581
rect 199 547 417 581
rect -417 -581 -199 -547
rect -109 -581 109 -547
rect 199 -581 417 -547
<< locali >>
rect -593 649 -497 683
rect 497 649 593 683
rect -593 587 -559 649
rect 559 587 593 649
rect -433 547 -417 581
rect -199 547 -183 581
rect -125 547 -109 581
rect 109 547 125 581
rect 183 547 199 581
rect 417 547 433 581
rect -479 488 -445 504
rect -479 -504 -445 -488
rect -171 488 -137 504
rect -171 -504 -137 -488
rect 137 488 171 504
rect 137 -504 171 -488
rect 445 488 479 504
rect 445 -504 479 -488
rect -433 -581 -417 -547
rect -199 -581 -183 -547
rect -125 -581 -109 -547
rect 109 -581 125 -547
rect 183 -581 199 -547
rect 417 -581 433 -547
rect -593 -649 -559 -587
rect 559 -649 593 -587
rect -593 -683 -497 -649
rect 497 -683 593 -649
<< viali >>
rect -417 547 -199 581
rect -109 547 109 581
rect 199 547 417 581
rect -479 -488 -445 488
rect -171 -488 -137 488
rect 137 -488 171 488
rect 445 -488 479 488
rect -417 -581 -199 -547
rect -109 -581 109 -547
rect 199 -581 417 -547
<< metal1 >>
rect -429 581 -187 587
rect -429 547 -417 581
rect -199 547 -187 581
rect -429 541 -187 547
rect -121 581 121 587
rect -121 547 -109 581
rect 109 547 121 581
rect -121 541 121 547
rect 187 581 429 587
rect 187 547 199 581
rect 417 547 429 581
rect 187 541 429 547
rect -485 488 -439 500
rect -485 -488 -479 488
rect -445 -488 -439 488
rect -485 -500 -439 -488
rect -177 488 -131 500
rect -177 -488 -171 488
rect -137 -488 -131 488
rect -177 -500 -131 -488
rect 131 488 177 500
rect 131 -488 137 488
rect 171 -488 177 488
rect 131 -500 177 -488
rect 439 488 485 500
rect 439 -488 445 488
rect 479 -488 485 488
rect 439 -500 485 -488
rect -429 -547 -187 -541
rect -429 -581 -417 -547
rect -199 -581 -187 -547
rect -429 -587 -187 -581
rect -121 -547 121 -541
rect -121 -581 -109 -547
rect 109 -581 121 -547
rect -121 -587 121 -581
rect 187 -547 429 -541
rect 187 -581 199 -547
rect 417 -581 429 -547
rect 187 -587 429 -581
<< properties >>
string FIXED_BBOX -576 -666 576 666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 1.25 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
