magic
tech sky130A
magscale 1 2
timestamp 1664842101
<< locali >>
rect -44 4828 14 4842
rect -44 2894 -32 4828
rect 2 2894 14 4828
rect 258 4808 274 4842
rect 310 4808 326 4842
rect 574 4808 590 4842
rect 626 4808 642 4842
rect 890 4808 906 4842
rect 942 4808 958 4842
rect 1206 4808 1222 4842
rect 1258 4808 1274 4842
rect 1522 4808 1538 4842
rect 1574 4808 1590 4842
rect 1838 4808 1854 4842
rect 1890 4808 1906 4842
rect 2154 4808 2170 4842
rect 2206 4808 2222 4842
rect 2470 4808 2486 4842
rect 2522 4808 2538 4842
rect 2786 4808 2802 4842
rect 2838 4808 2854 4842
rect 3102 4808 3118 4842
rect 3154 4808 3170 4842
rect 3418 4808 3434 4842
rect 3470 4808 3486 4842
rect 3734 4808 3750 4842
rect 3786 4808 3802 4842
rect 4050 4808 4066 4842
rect 4102 4808 4118 4842
rect 4366 4808 4382 4842
rect 4418 4808 4434 4842
rect 4682 4808 4698 4842
rect 4734 4808 4750 4842
rect 4998 4808 5014 4842
rect 5050 4808 5066 4842
rect 5314 4808 5330 4842
rect 5366 4808 5382 4842
rect 5630 4808 5646 4842
rect 5682 4808 5698 4842
rect 5946 4808 5962 4842
rect 5998 4808 6014 4842
rect 6262 4808 6278 4842
rect 6314 4808 6330 4842
rect 6578 4808 6594 4842
rect 6630 4808 6646 4842
rect 6894 4808 6910 4842
rect 6946 4808 6962 4842
rect 7210 4808 7226 4842
rect 7262 4808 7278 4842
rect 7526 4808 7542 4842
rect 7578 4808 7594 4842
rect 7842 4808 7858 4842
rect 7894 4808 7910 4842
rect 8158 4808 8174 4842
rect 8210 4808 8226 4842
rect 8474 4808 8490 4842
rect 8526 4808 8542 4842
rect 8790 4808 8806 4842
rect 8842 4808 8858 4842
rect 9106 4808 9122 4842
rect 9158 4808 9174 4842
rect 9422 4808 9438 4842
rect 9474 4808 9490 4842
rect 9738 4808 9754 4842
rect 9790 4808 9806 4842
rect 10054 4808 10070 4842
rect 10106 4808 10122 4842
rect 10370 4808 10386 4842
rect 10422 4808 10438 4842
rect 10686 4808 10702 4842
rect 10738 4808 10754 4842
rect 11002 4808 11018 4842
rect 11054 4808 11070 4842
rect 11318 4808 11334 4842
rect 11370 4808 11386 4842
rect 11634 4808 11650 4842
rect 11686 4808 11702 4842
rect 11950 4808 11966 4842
rect 12002 4808 12018 4842
rect 12266 4808 12282 4842
rect 12318 4808 12334 4842
rect 12582 4808 12598 4842
rect 12634 4808 12650 4842
rect 12892 4828 12950 4842
rect -44 2854 14 2894
rect 12892 2894 12904 4828
rect 12938 2894 12950 4828
rect 12892 2854 12950 2894
rect -44 1932 14 1972
rect -44 -6 -32 1932
rect 2 -6 14 1932
rect 12892 1932 12950 1972
rect -44 -18 14 -6
rect 268 -18 274 16
rect 310 -18 316 16
rect 574 -18 590 16
rect 626 -18 642 16
rect 890 -18 906 16
rect 942 -18 958 16
rect 1206 -18 1222 16
rect 1258 -18 1274 16
rect 1522 -18 1538 16
rect 1574 -18 1590 16
rect 1838 -18 1854 16
rect 1890 -18 1906 16
rect 2154 -18 2170 16
rect 2206 -18 2222 16
rect 2470 -18 2486 16
rect 2522 -18 2538 16
rect 2786 -18 2802 16
rect 2838 -18 2854 16
rect 3102 -18 3118 16
rect 3154 -18 3170 16
rect 3418 -18 3434 16
rect 3470 -18 3486 16
rect 3734 -18 3750 16
rect 3786 -18 3802 16
rect 4050 -18 4066 16
rect 4102 -18 4118 16
rect 4366 -18 4382 16
rect 4418 -18 4434 16
rect 4682 -18 4698 16
rect 4734 -18 4750 16
rect 4998 -18 5014 16
rect 5050 -18 5066 16
rect 5314 -18 5330 16
rect 5366 -18 5382 16
rect 5630 -18 5646 16
rect 5682 -18 5698 16
rect 5946 -18 5962 16
rect 5998 -18 6014 16
rect 6262 -18 6278 16
rect 6314 -18 6330 16
rect 6578 -18 6594 16
rect 6630 -18 6646 16
rect 6894 -18 6910 16
rect 6946 -18 6962 16
rect 7210 -18 7226 16
rect 7262 -18 7278 16
rect 7526 -18 7542 16
rect 7578 -18 7594 16
rect 7842 -18 7858 16
rect 7894 -18 7910 16
rect 8158 -18 8174 16
rect 8210 -18 8226 16
rect 8474 -18 8490 16
rect 8526 -18 8542 16
rect 8790 -18 8806 16
rect 8842 -18 8858 16
rect 9106 -18 9122 16
rect 9158 -18 9174 16
rect 9422 -18 9438 16
rect 9474 -18 9490 16
rect 9738 -18 9754 16
rect 9790 -18 9806 16
rect 10054 -18 10070 16
rect 10106 -18 10122 16
rect 10370 -18 10386 16
rect 10422 -18 10438 16
rect 10686 -18 10702 16
rect 10738 -18 10754 16
rect 11002 -18 11018 16
rect 11054 -18 11070 16
rect 11318 -18 11334 16
rect 11370 -18 11386 16
rect 11634 -18 11650 16
rect 11686 -18 11702 16
rect 11950 -18 11966 16
rect 12002 -18 12018 16
rect 12266 -18 12282 16
rect 12318 -18 12334 16
rect 12582 -18 12598 16
rect 12634 -18 12650 16
rect 12892 -6 12904 1932
rect 12938 -6 12950 1932
rect 12892 -18 12950 -6
<< viali >>
rect -32 2894 2 4828
rect 274 4808 310 4842
rect 590 4808 626 4842
rect 906 4808 942 4842
rect 1222 4808 1258 4842
rect 1538 4808 1574 4842
rect 1854 4808 1890 4842
rect 2170 4808 2206 4842
rect 2486 4808 2522 4842
rect 2802 4808 2838 4842
rect 3118 4808 3154 4842
rect 3434 4808 3470 4842
rect 3750 4808 3786 4842
rect 4066 4808 4102 4842
rect 4382 4808 4418 4842
rect 4698 4808 4734 4842
rect 5014 4808 5050 4842
rect 5330 4808 5366 4842
rect 5646 4808 5682 4842
rect 5962 4808 5998 4842
rect 6278 4808 6314 4842
rect 6594 4808 6630 4842
rect 6910 4808 6946 4842
rect 7226 4808 7262 4842
rect 7542 4808 7578 4842
rect 7858 4808 7894 4842
rect 8174 4808 8210 4842
rect 8490 4808 8526 4842
rect 8806 4808 8842 4842
rect 9122 4808 9158 4842
rect 9438 4808 9474 4842
rect 9754 4808 9790 4842
rect 10070 4808 10106 4842
rect 10386 4808 10422 4842
rect 10702 4808 10738 4842
rect 11018 4808 11054 4842
rect 11334 4808 11370 4842
rect 11650 4808 11686 4842
rect 11966 4808 12002 4842
rect 12282 4808 12318 4842
rect 12598 4808 12634 4842
rect 12904 2894 12938 4828
rect -32 -6 2 1932
rect 274 -18 310 16
rect 590 -18 626 16
rect 906 -18 942 16
rect 1222 -18 1258 16
rect 1538 -18 1574 16
rect 1854 -18 1890 16
rect 2170 -18 2206 16
rect 2486 -18 2522 16
rect 2802 -18 2838 16
rect 3118 -18 3154 16
rect 3434 -18 3470 16
rect 3750 -18 3786 16
rect 4066 -18 4102 16
rect 4382 -18 4418 16
rect 4698 -18 4734 16
rect 5014 -18 5050 16
rect 5330 -18 5366 16
rect 5646 -18 5682 16
rect 5962 -18 5998 16
rect 6278 -18 6314 16
rect 6594 -18 6630 16
rect 6910 -18 6946 16
rect 7226 -18 7262 16
rect 7542 -18 7578 16
rect 7858 -18 7894 16
rect 8174 -18 8210 16
rect 8490 -18 8526 16
rect 8806 -18 8842 16
rect 9122 -18 9158 16
rect 9438 -18 9474 16
rect 9754 -18 9790 16
rect 10070 -18 10106 16
rect 10386 -18 10422 16
rect 10702 -18 10738 16
rect 11018 -18 11054 16
rect 11334 -18 11370 16
rect 11650 -18 11686 16
rect 11966 -18 12002 16
rect 12282 -18 12318 16
rect 12598 -18 12634 16
rect 12904 -6 12938 1932
<< metal1 >>
rect 254 4852 330 4858
rect 254 4842 260 4852
rect 324 4842 330 4852
rect 570 4852 646 4858
rect 570 4842 576 4852
rect 640 4842 646 4852
rect 886 4852 962 4858
rect 886 4842 892 4852
rect 956 4842 962 4852
rect 1202 4852 1278 4858
rect 1202 4842 1208 4852
rect 1272 4842 1278 4852
rect 1518 4852 1594 4858
rect 1518 4842 1524 4852
rect 1588 4842 1594 4852
rect 1834 4852 1910 4858
rect 1834 4842 1840 4852
rect 1904 4842 1910 4852
rect 2150 4852 2226 4858
rect 2150 4842 2156 4852
rect 2220 4842 2226 4852
rect 2466 4852 2542 4858
rect 2466 4842 2472 4852
rect 2536 4842 2542 4852
rect 2782 4852 2858 4858
rect 2782 4842 2788 4852
rect 2852 4842 2858 4852
rect 3098 4852 3174 4858
rect 3098 4842 3104 4852
rect 3168 4842 3174 4852
rect 3414 4852 3490 4858
rect 3414 4842 3420 4852
rect 3484 4842 3490 4852
rect 3730 4852 3806 4858
rect 3730 4842 3736 4852
rect 3800 4842 3806 4852
rect 4046 4852 4122 4858
rect 4046 4842 4052 4852
rect 4116 4842 4122 4852
rect 4362 4852 4438 4858
rect 4362 4842 4368 4852
rect 4432 4842 4438 4852
rect 4678 4852 4754 4858
rect 4678 4842 4684 4852
rect 4748 4842 4754 4852
rect 4994 4852 5070 4858
rect 4994 4842 5000 4852
rect 5064 4842 5070 4852
rect 5310 4852 5386 4858
rect 5310 4842 5316 4852
rect 5380 4842 5386 4852
rect 5626 4852 5702 4858
rect 5626 4842 5632 4852
rect 5696 4842 5702 4852
rect 5942 4852 6018 4858
rect 5942 4842 5948 4852
rect 6012 4842 6018 4852
rect 6258 4852 6334 4858
rect 6258 4842 6264 4852
rect 6328 4842 6334 4852
rect 6574 4852 6650 4858
rect 6574 4842 6580 4852
rect 6644 4842 6650 4852
rect 6890 4852 6966 4858
rect 6890 4842 6896 4852
rect 6960 4842 6966 4852
rect 7206 4852 7282 4858
rect 7206 4842 7212 4852
rect 7276 4842 7282 4852
rect 7522 4852 7598 4858
rect 7522 4842 7528 4852
rect 7592 4842 7598 4852
rect 7838 4852 7914 4858
rect 7838 4842 7844 4852
rect 7908 4842 7914 4852
rect 8154 4852 8230 4858
rect 8154 4842 8160 4852
rect 8224 4842 8230 4852
rect 8470 4852 8546 4858
rect 8470 4842 8476 4852
rect 8540 4842 8546 4852
rect 8786 4852 8862 4858
rect 8786 4842 8792 4852
rect 8856 4842 8862 4852
rect 9102 4852 9178 4858
rect 9102 4842 9108 4852
rect 9172 4842 9178 4852
rect 9418 4852 9494 4858
rect 9418 4842 9424 4852
rect 9488 4842 9494 4852
rect 9734 4852 9810 4858
rect 9734 4842 9740 4852
rect 9804 4842 9810 4852
rect 10050 4852 10126 4858
rect 10050 4842 10056 4852
rect 10120 4842 10126 4852
rect 10366 4852 10442 4858
rect 10366 4842 10372 4852
rect 10436 4842 10442 4852
rect 10682 4852 10758 4858
rect 10682 4842 10688 4852
rect 10752 4842 10758 4852
rect 10998 4852 11074 4858
rect 10998 4842 11004 4852
rect 11068 4842 11074 4852
rect 11314 4852 11390 4858
rect 11314 4842 11320 4852
rect 11384 4842 11390 4852
rect 11630 4852 11706 4858
rect 11630 4842 11636 4852
rect 11700 4842 11706 4852
rect 11946 4852 12022 4858
rect 11946 4842 11952 4852
rect 12016 4842 12022 4852
rect 12262 4852 12338 4858
rect 12262 4842 12268 4852
rect 12332 4842 12338 4852
rect 12578 4852 12654 4858
rect 12578 4842 12584 4852
rect 12648 4842 12654 4852
rect -44 4828 260 4842
rect -44 2894 -32 4828
rect 2 4808 260 4828
rect 324 4808 576 4842
rect 640 4808 892 4842
rect 956 4808 1208 4842
rect 1272 4808 1524 4842
rect 1588 4808 1840 4842
rect 1904 4808 2156 4842
rect 2220 4808 2472 4842
rect 2536 4808 2788 4842
rect 2852 4808 3104 4842
rect 3168 4808 3420 4842
rect 3484 4808 3736 4842
rect 3800 4808 4052 4842
rect 4116 4808 4368 4842
rect 4432 4808 4684 4842
rect 4748 4808 5000 4842
rect 5064 4808 5316 4842
rect 5380 4808 5632 4842
rect 5696 4808 5948 4842
rect 6012 4808 6264 4842
rect 6328 4808 6580 4842
rect 6644 4808 6896 4842
rect 6960 4808 7212 4842
rect 7276 4808 7528 4842
rect 7592 4808 7844 4842
rect 7908 4808 8160 4842
rect 8224 4808 8476 4842
rect 8540 4808 8792 4842
rect 8856 4808 9108 4842
rect 9172 4808 9424 4842
rect 9488 4808 9740 4842
rect 9804 4808 10056 4842
rect 10120 4808 10372 4842
rect 10436 4808 10688 4842
rect 10752 4808 11004 4842
rect 11068 4808 11320 4842
rect 11384 4808 11636 4842
rect 11700 4808 11952 4842
rect 12016 4808 12268 4842
rect 12332 4808 12584 4842
rect 12648 4828 12950 4842
rect 12648 4808 12904 4828
rect 2 2894 14 4808
rect 254 4798 260 4808
rect 324 4798 330 4808
rect 254 4792 330 4798
rect 570 4798 576 4808
rect 640 4798 646 4808
rect 570 4792 646 4798
rect 886 4798 892 4808
rect 956 4798 962 4808
rect 886 4792 962 4798
rect 1202 4798 1208 4808
rect 1272 4798 1278 4808
rect 1202 4792 1278 4798
rect 1518 4798 1524 4808
rect 1588 4798 1594 4808
rect 1518 4792 1594 4798
rect 1834 4798 1840 4808
rect 1904 4798 1910 4808
rect 1834 4792 1910 4798
rect 2150 4798 2156 4808
rect 2220 4798 2226 4808
rect 2150 4792 2226 4798
rect 2466 4798 2472 4808
rect 2536 4798 2542 4808
rect 2466 4792 2542 4798
rect 2782 4798 2788 4808
rect 2852 4798 2858 4808
rect 2782 4792 2858 4798
rect 3098 4798 3104 4808
rect 3168 4798 3174 4808
rect 3098 4792 3174 4798
rect 3414 4798 3420 4808
rect 3484 4798 3490 4808
rect 3414 4792 3490 4798
rect 3730 4798 3736 4808
rect 3800 4798 3806 4808
rect 3730 4792 3806 4798
rect 4046 4798 4052 4808
rect 4116 4798 4122 4808
rect 4046 4792 4122 4798
rect 4362 4798 4368 4808
rect 4432 4798 4438 4808
rect 4362 4792 4438 4798
rect 4678 4798 4684 4808
rect 4748 4798 4754 4808
rect 4678 4792 4754 4798
rect 4994 4798 5000 4808
rect 5064 4798 5070 4808
rect 4994 4792 5070 4798
rect 5310 4798 5316 4808
rect 5380 4798 5386 4808
rect 5310 4792 5386 4798
rect 5626 4798 5632 4808
rect 5696 4798 5702 4808
rect 5626 4792 5702 4798
rect 5942 4798 5948 4808
rect 6012 4798 6018 4808
rect 5942 4792 6018 4798
rect 6258 4798 6264 4808
rect 6328 4798 6334 4808
rect 6258 4792 6334 4798
rect 6574 4798 6580 4808
rect 6644 4798 6650 4808
rect 6574 4792 6650 4798
rect 6890 4798 6896 4808
rect 6960 4798 6966 4808
rect 6890 4792 6966 4798
rect 7206 4798 7212 4808
rect 7276 4798 7282 4808
rect 7206 4792 7282 4798
rect 7522 4798 7528 4808
rect 7592 4798 7598 4808
rect 7522 4792 7598 4798
rect 7838 4798 7844 4808
rect 7908 4798 7914 4808
rect 7838 4792 7914 4798
rect 8154 4798 8160 4808
rect 8224 4798 8230 4808
rect 8154 4792 8230 4798
rect 8470 4798 8476 4808
rect 8540 4798 8546 4808
rect 8470 4792 8546 4798
rect 8786 4798 8792 4808
rect 8856 4798 8862 4808
rect 8786 4792 8862 4798
rect 9102 4798 9108 4808
rect 9172 4798 9178 4808
rect 9102 4792 9178 4798
rect 9418 4798 9424 4808
rect 9488 4798 9494 4808
rect 9418 4792 9494 4798
rect 9734 4798 9740 4808
rect 9804 4798 9810 4808
rect 9734 4792 9810 4798
rect 10050 4798 10056 4808
rect 10120 4798 10126 4808
rect 10050 4792 10126 4798
rect 10366 4798 10372 4808
rect 10436 4798 10442 4808
rect 10366 4792 10442 4798
rect 10682 4798 10688 4808
rect 10752 4798 10758 4808
rect 10682 4792 10758 4798
rect 10998 4798 11004 4808
rect 11068 4798 11074 4808
rect 10998 4792 11074 4798
rect 11314 4798 11320 4808
rect 11384 4798 11390 4808
rect 11314 4792 11390 4798
rect 11630 4798 11636 4808
rect 11700 4798 11706 4808
rect 11630 4792 11706 4798
rect 11946 4798 11952 4808
rect 12016 4798 12022 4808
rect 11946 4792 12022 4798
rect 12262 4798 12268 4808
rect 12332 4798 12338 4808
rect 12262 4792 12338 4798
rect 12578 4798 12584 4808
rect 12648 4798 12654 4808
rect 12578 4792 12654 4798
rect -44 2854 14 2894
rect 42 4664 12864 4711
rect 42 3800 76 4664
rect 104 4622 168 4628
rect 269 4626 315 4632
rect 427 4628 473 4632
rect 104 3844 110 4622
rect 162 3844 168 4622
rect 104 3838 168 3844
rect 262 4622 326 4626
rect 262 3840 268 4622
rect 320 3840 326 4622
rect 262 3836 326 3840
rect 420 4622 484 4628
rect 585 4626 631 4632
rect 743 4628 789 4632
rect 420 3844 426 4622
rect 478 3844 484 4622
rect 420 3838 484 3844
rect 578 4622 642 4626
rect 578 3840 584 4622
rect 636 3840 642 4622
rect 269 3832 315 3836
rect 427 3832 473 3838
rect 578 3836 642 3840
rect 736 4622 800 4628
rect 901 4626 947 4632
rect 1059 4628 1105 4632
rect 736 3844 742 4622
rect 794 3844 800 4622
rect 736 3838 800 3844
rect 894 4622 958 4626
rect 894 3840 900 4622
rect 952 3840 958 4622
rect 585 3832 631 3836
rect 743 3832 789 3838
rect 894 3836 958 3840
rect 1052 4622 1116 4628
rect 1217 4626 1263 4632
rect 1375 4628 1421 4632
rect 1052 3844 1058 4622
rect 1110 3844 1116 4622
rect 1052 3838 1116 3844
rect 1210 4622 1274 4626
rect 1210 3840 1216 4622
rect 1268 3840 1274 4622
rect 901 3832 947 3836
rect 1059 3832 1105 3838
rect 1210 3836 1274 3840
rect 1368 4622 1432 4628
rect 1533 4626 1579 4632
rect 1691 4628 1737 4632
rect 1368 3844 1374 4622
rect 1426 3844 1432 4622
rect 1368 3838 1432 3844
rect 1526 4622 1590 4626
rect 1526 3840 1532 4622
rect 1584 3840 1590 4622
rect 1217 3832 1263 3836
rect 1375 3832 1421 3838
rect 1526 3836 1590 3840
rect 1684 4622 1748 4628
rect 1849 4626 1895 4632
rect 2007 4628 2053 4632
rect 1684 3844 1690 4622
rect 1742 3844 1748 4622
rect 1684 3838 1748 3844
rect 1842 4622 1906 4626
rect 1842 3840 1848 4622
rect 1900 3840 1906 4622
rect 1533 3832 1579 3836
rect 1691 3832 1737 3838
rect 1842 3836 1906 3840
rect 2000 4622 2064 4628
rect 2165 4626 2211 4632
rect 2323 4628 2369 4632
rect 2000 3844 2006 4622
rect 2058 3844 2064 4622
rect 2000 3838 2064 3844
rect 2158 4622 2222 4626
rect 2158 3840 2164 4622
rect 2216 3840 2222 4622
rect 1849 3832 1895 3836
rect 2007 3832 2053 3838
rect 2158 3836 2222 3840
rect 2316 4622 2380 4628
rect 2481 4626 2527 4632
rect 2639 4628 2685 4632
rect 2316 3844 2322 4622
rect 2374 3844 2380 4622
rect 2316 3838 2380 3844
rect 2474 4622 2538 4626
rect 2474 3840 2480 4622
rect 2532 3840 2538 4622
rect 2165 3832 2211 3836
rect 2323 3832 2369 3838
rect 2474 3836 2538 3840
rect 2632 4622 2696 4628
rect 2797 4626 2843 4632
rect 2955 4628 3001 4632
rect 2632 3844 2638 4622
rect 2690 3844 2696 4622
rect 2632 3838 2696 3844
rect 2790 4622 2854 4626
rect 2790 3840 2796 4622
rect 2848 3840 2854 4622
rect 2481 3832 2527 3836
rect 2639 3832 2685 3838
rect 2790 3836 2854 3840
rect 2948 4622 3012 4628
rect 3113 4626 3159 4632
rect 3271 4628 3317 4632
rect 2948 3844 2954 4622
rect 3006 3844 3012 4622
rect 2948 3838 3012 3844
rect 3106 4622 3170 4626
rect 3106 3840 3112 4622
rect 3164 3840 3170 4622
rect 2797 3832 2843 3836
rect 2955 3832 3001 3838
rect 3106 3836 3170 3840
rect 3264 4622 3328 4628
rect 3429 4626 3475 4632
rect 3587 4628 3633 4632
rect 3264 3844 3270 4622
rect 3322 3844 3328 4622
rect 3264 3838 3328 3844
rect 3422 4622 3486 4626
rect 3422 3840 3428 4622
rect 3480 3840 3486 4622
rect 3113 3832 3159 3836
rect 3271 3832 3317 3838
rect 3422 3836 3486 3840
rect 3580 4622 3644 4628
rect 3745 4626 3791 4632
rect 3903 4628 3949 4632
rect 3580 3844 3586 4622
rect 3638 3844 3644 4622
rect 3580 3838 3644 3844
rect 3738 4622 3802 4626
rect 3738 3840 3744 4622
rect 3796 3840 3802 4622
rect 3429 3832 3475 3836
rect 3587 3832 3633 3838
rect 3738 3836 3802 3840
rect 3896 4622 3960 4628
rect 4061 4626 4107 4632
rect 4219 4628 4265 4632
rect 3896 3844 3902 4622
rect 3954 3844 3960 4622
rect 3896 3838 3960 3844
rect 4054 4622 4118 4626
rect 4054 3840 4060 4622
rect 4112 3840 4118 4622
rect 3745 3832 3791 3836
rect 3903 3832 3949 3838
rect 4054 3836 4118 3840
rect 4212 4622 4276 4628
rect 4377 4626 4423 4632
rect 4535 4628 4581 4632
rect 4212 3844 4218 4622
rect 4270 3844 4276 4622
rect 4212 3838 4276 3844
rect 4370 4622 4434 4626
rect 4370 3840 4376 4622
rect 4428 3840 4434 4622
rect 4061 3832 4107 3836
rect 4219 3832 4265 3838
rect 4370 3836 4434 3840
rect 4528 4622 4592 4628
rect 4693 4626 4739 4632
rect 4851 4628 4897 4632
rect 4528 3844 4534 4622
rect 4586 3844 4592 4622
rect 4528 3838 4592 3844
rect 4686 4622 4750 4626
rect 4686 3840 4692 4622
rect 4744 3840 4750 4622
rect 4377 3832 4423 3836
rect 4535 3832 4581 3838
rect 4686 3836 4750 3840
rect 4844 4622 4908 4628
rect 5009 4626 5055 4632
rect 5167 4628 5213 4632
rect 4844 3844 4850 4622
rect 4902 3844 4908 4622
rect 4844 3838 4908 3844
rect 5002 4622 5066 4626
rect 5002 3840 5008 4622
rect 5060 3840 5066 4622
rect 4693 3832 4739 3836
rect 4851 3832 4897 3838
rect 5002 3836 5066 3840
rect 5160 4622 5224 4628
rect 5325 4626 5371 4632
rect 5483 4628 5529 4632
rect 5160 3844 5166 4622
rect 5218 3844 5224 4622
rect 5160 3838 5224 3844
rect 5318 4622 5382 4626
rect 5318 3840 5324 4622
rect 5376 3840 5382 4622
rect 5009 3832 5055 3836
rect 5167 3832 5213 3838
rect 5318 3836 5382 3840
rect 5476 4622 5540 4628
rect 5641 4626 5687 4632
rect 5799 4628 5845 4632
rect 5476 3844 5482 4622
rect 5534 3844 5540 4622
rect 5476 3838 5540 3844
rect 5634 4622 5698 4626
rect 5634 3840 5640 4622
rect 5692 3840 5698 4622
rect 5325 3832 5371 3836
rect 5483 3832 5529 3838
rect 5634 3836 5698 3840
rect 5792 4622 5856 4628
rect 5957 4626 6003 4632
rect 6115 4628 6161 4632
rect 5792 3844 5798 4622
rect 5850 3844 5856 4622
rect 5792 3838 5856 3844
rect 5950 4622 6014 4626
rect 5950 3840 5956 4622
rect 6008 3840 6014 4622
rect 5641 3832 5687 3836
rect 5799 3832 5845 3838
rect 5950 3836 6014 3840
rect 6108 4622 6172 4628
rect 6273 4626 6319 4632
rect 6431 4628 6477 4632
rect 6108 3844 6114 4622
rect 6166 3844 6172 4622
rect 6108 3838 6172 3844
rect 6266 4622 6330 4626
rect 6266 3840 6272 4622
rect 6324 3840 6330 4622
rect 5957 3832 6003 3836
rect 6115 3832 6161 3838
rect 6266 3836 6330 3840
rect 6424 4622 6488 4628
rect 6589 4626 6635 4632
rect 6747 4628 6793 4632
rect 6424 3844 6430 4622
rect 6482 3844 6488 4622
rect 6424 3838 6488 3844
rect 6582 4622 6646 4626
rect 6582 3840 6588 4622
rect 6640 3840 6646 4622
rect 6273 3832 6319 3836
rect 6431 3832 6477 3838
rect 6582 3836 6646 3840
rect 6740 4622 6804 4628
rect 6905 4626 6951 4632
rect 7063 4628 7109 4632
rect 6740 3844 6746 4622
rect 6798 3844 6804 4622
rect 6740 3838 6804 3844
rect 6898 4622 6962 4626
rect 6898 3840 6904 4622
rect 6956 3840 6962 4622
rect 6589 3832 6635 3836
rect 6747 3832 6793 3838
rect 6898 3836 6962 3840
rect 7056 4622 7120 4628
rect 7221 4626 7267 4632
rect 7379 4628 7425 4632
rect 7056 3844 7062 4622
rect 7114 3844 7120 4622
rect 7056 3838 7120 3844
rect 7214 4622 7278 4626
rect 7214 3840 7220 4622
rect 7272 3840 7278 4622
rect 6905 3832 6951 3836
rect 7063 3832 7109 3838
rect 7214 3836 7278 3840
rect 7372 4622 7436 4628
rect 7537 4626 7583 4632
rect 7695 4628 7741 4632
rect 7372 3844 7378 4622
rect 7430 3844 7436 4622
rect 7372 3838 7436 3844
rect 7530 4622 7594 4626
rect 7530 3840 7536 4622
rect 7588 3840 7594 4622
rect 7221 3832 7267 3836
rect 7379 3832 7425 3838
rect 7530 3836 7594 3840
rect 7688 4622 7752 4628
rect 7853 4626 7899 4632
rect 8011 4628 8057 4632
rect 7688 3844 7694 4622
rect 7746 3844 7752 4622
rect 7688 3838 7752 3844
rect 7846 4622 7910 4626
rect 7846 3840 7852 4622
rect 7904 3840 7910 4622
rect 7537 3832 7583 3836
rect 7695 3832 7741 3838
rect 7846 3836 7910 3840
rect 8004 4622 8068 4628
rect 8169 4626 8215 4632
rect 8327 4628 8373 4632
rect 8004 3844 8010 4622
rect 8062 3844 8068 4622
rect 8004 3838 8068 3844
rect 8162 4622 8226 4626
rect 8162 3840 8168 4622
rect 8220 3840 8226 4622
rect 7853 3832 7899 3836
rect 8011 3832 8057 3838
rect 8162 3836 8226 3840
rect 8320 4622 8384 4628
rect 8485 4626 8531 4632
rect 8643 4628 8689 4632
rect 8320 3844 8326 4622
rect 8378 3844 8384 4622
rect 8320 3838 8384 3844
rect 8478 4622 8542 4626
rect 8478 3840 8484 4622
rect 8536 3840 8542 4622
rect 8169 3832 8215 3836
rect 8327 3832 8373 3838
rect 8478 3836 8542 3840
rect 8636 4622 8700 4628
rect 8801 4626 8847 4632
rect 8959 4628 9005 4632
rect 8636 3844 8642 4622
rect 8694 3844 8700 4622
rect 8636 3838 8700 3844
rect 8794 4622 8858 4626
rect 8794 3840 8800 4622
rect 8852 3840 8858 4622
rect 8485 3832 8531 3836
rect 8643 3832 8689 3838
rect 8794 3836 8858 3840
rect 8952 4622 9016 4628
rect 9117 4626 9163 4632
rect 9275 4628 9321 4632
rect 8952 3844 8958 4622
rect 9010 3844 9016 4622
rect 8952 3838 9016 3844
rect 9110 4622 9174 4626
rect 9110 3840 9116 4622
rect 9168 3840 9174 4622
rect 8801 3832 8847 3836
rect 8959 3832 9005 3838
rect 9110 3836 9174 3840
rect 9268 4622 9332 4628
rect 9433 4626 9479 4632
rect 9591 4628 9637 4632
rect 9268 3844 9274 4622
rect 9326 3844 9332 4622
rect 9268 3838 9332 3844
rect 9426 4622 9490 4626
rect 9426 3840 9432 4622
rect 9484 3840 9490 4622
rect 9117 3832 9163 3836
rect 9275 3832 9321 3838
rect 9426 3836 9490 3840
rect 9584 4622 9648 4628
rect 9749 4626 9795 4632
rect 9907 4628 9953 4632
rect 9584 3844 9590 4622
rect 9642 3844 9648 4622
rect 9584 3838 9648 3844
rect 9742 4622 9806 4626
rect 9742 3840 9748 4622
rect 9800 3840 9806 4622
rect 9433 3832 9479 3836
rect 9591 3832 9637 3838
rect 9742 3836 9806 3840
rect 9900 4622 9964 4628
rect 10065 4626 10111 4632
rect 10223 4628 10269 4632
rect 9900 3844 9906 4622
rect 9958 3844 9964 4622
rect 9900 3838 9964 3844
rect 10058 4622 10122 4626
rect 10058 3840 10064 4622
rect 10116 3840 10122 4622
rect 9749 3832 9795 3836
rect 9907 3832 9953 3838
rect 10058 3836 10122 3840
rect 10216 4622 10280 4628
rect 10381 4626 10427 4632
rect 10539 4628 10585 4632
rect 10216 3844 10222 4622
rect 10274 3844 10280 4622
rect 10216 3838 10280 3844
rect 10374 4622 10438 4626
rect 10374 3840 10380 4622
rect 10432 3840 10438 4622
rect 10065 3832 10111 3836
rect 10223 3832 10269 3838
rect 10374 3836 10438 3840
rect 10532 4622 10596 4628
rect 10697 4626 10743 4632
rect 10855 4628 10901 4632
rect 10532 3844 10538 4622
rect 10590 3844 10596 4622
rect 10532 3838 10596 3844
rect 10690 4622 10754 4626
rect 10690 3840 10696 4622
rect 10748 3840 10754 4622
rect 10381 3832 10427 3836
rect 10539 3832 10585 3838
rect 10690 3836 10754 3840
rect 10848 4622 10912 4628
rect 11013 4626 11059 4632
rect 11171 4628 11217 4632
rect 10848 3844 10854 4622
rect 10906 3844 10912 4622
rect 10848 3838 10912 3844
rect 11006 4622 11070 4626
rect 11006 3840 11012 4622
rect 11064 3840 11070 4622
rect 10697 3832 10743 3836
rect 10855 3832 10901 3838
rect 11006 3836 11070 3840
rect 11164 4622 11228 4628
rect 11329 4626 11375 4632
rect 11487 4628 11533 4632
rect 11164 3844 11170 4622
rect 11222 3844 11228 4622
rect 11164 3838 11228 3844
rect 11322 4622 11386 4626
rect 11322 3840 11328 4622
rect 11380 3840 11386 4622
rect 11013 3832 11059 3836
rect 11171 3832 11217 3838
rect 11322 3836 11386 3840
rect 11480 4622 11544 4628
rect 11645 4626 11691 4632
rect 11803 4628 11849 4632
rect 11480 3844 11486 4622
rect 11538 3844 11544 4622
rect 11480 3838 11544 3844
rect 11638 4622 11702 4626
rect 11638 3840 11644 4622
rect 11696 3840 11702 4622
rect 11329 3832 11375 3836
rect 11487 3832 11533 3838
rect 11638 3836 11702 3840
rect 11796 4622 11860 4628
rect 11961 4626 12007 4632
rect 12119 4628 12165 4632
rect 11796 3844 11802 4622
rect 11854 3844 11860 4622
rect 11796 3838 11860 3844
rect 11954 4622 12018 4626
rect 11954 3840 11960 4622
rect 12012 3840 12018 4622
rect 11645 3832 11691 3836
rect 11803 3832 11849 3838
rect 11954 3836 12018 3840
rect 12112 4622 12176 4628
rect 12277 4626 12323 4632
rect 12435 4628 12481 4632
rect 12112 3844 12118 4622
rect 12170 3844 12176 4622
rect 12112 3838 12176 3844
rect 12270 4622 12334 4626
rect 12270 3840 12276 4622
rect 12328 3840 12334 4622
rect 11961 3832 12007 3836
rect 12119 3832 12165 3838
rect 12270 3836 12334 3840
rect 12428 4622 12492 4628
rect 12593 4626 12639 4632
rect 12745 4628 12791 4632
rect 12428 3844 12434 4622
rect 12486 3844 12492 4622
rect 12428 3838 12492 3844
rect 12586 4622 12650 4626
rect 12586 3840 12592 4622
rect 12644 3840 12650 4622
rect 12277 3832 12323 3836
rect 12435 3832 12481 3838
rect 12586 3836 12650 3840
rect 12738 4622 12802 4628
rect 12738 3844 12744 4622
rect 12796 3844 12802 4622
rect 12738 3838 12802 3844
rect 12593 3832 12639 3836
rect 12745 3832 12791 3838
rect 12830 3800 12864 4664
rect 42 3754 12864 3800
rect 42 2890 76 3754
rect 104 3714 168 3718
rect 269 3716 315 3722
rect 427 3718 473 3722
rect 104 2932 110 3714
rect 162 2932 168 3714
rect 104 2928 168 2932
rect 262 3712 326 3716
rect 262 2930 268 3712
rect 320 2930 326 3712
rect 262 2926 326 2930
rect 420 3714 484 3718
rect 585 3716 631 3722
rect 743 3718 789 3722
rect 420 2932 426 3714
rect 478 2932 484 3714
rect 420 2928 484 2932
rect 578 3712 642 3716
rect 578 2930 584 3712
rect 636 2930 642 3712
rect 269 2922 315 2926
rect 427 2922 473 2928
rect 578 2926 642 2930
rect 736 3714 800 3718
rect 901 3716 947 3722
rect 1059 3718 1105 3722
rect 736 2932 742 3714
rect 794 2932 800 3714
rect 736 2928 800 2932
rect 894 3712 958 3716
rect 894 2930 900 3712
rect 952 2930 958 3712
rect 585 2922 631 2926
rect 743 2922 789 2928
rect 894 2926 958 2930
rect 1052 3714 1116 3718
rect 1217 3716 1263 3722
rect 1375 3718 1421 3722
rect 1052 2932 1058 3714
rect 1110 2932 1116 3714
rect 1052 2928 1116 2932
rect 1210 3712 1274 3716
rect 1210 2930 1216 3712
rect 1268 2930 1274 3712
rect 901 2922 947 2926
rect 1059 2922 1105 2928
rect 1210 2926 1274 2930
rect 1368 3714 1432 3718
rect 1533 3716 1579 3722
rect 1691 3718 1737 3722
rect 1368 2932 1374 3714
rect 1426 2932 1432 3714
rect 1368 2928 1432 2932
rect 1526 3712 1590 3716
rect 1526 2930 1532 3712
rect 1584 2930 1590 3712
rect 1217 2922 1263 2926
rect 1375 2922 1421 2928
rect 1526 2926 1590 2930
rect 1684 3714 1748 3718
rect 1849 3716 1895 3722
rect 2007 3718 2053 3722
rect 1684 2932 1690 3714
rect 1742 2932 1748 3714
rect 1684 2928 1748 2932
rect 1842 3712 1906 3716
rect 1842 2930 1848 3712
rect 1900 2930 1906 3712
rect 1533 2922 1579 2926
rect 1691 2922 1737 2928
rect 1842 2926 1906 2930
rect 2000 3714 2064 3718
rect 2165 3716 2211 3722
rect 2323 3718 2369 3722
rect 2000 2932 2006 3714
rect 2058 2932 2064 3714
rect 2000 2928 2064 2932
rect 2158 3712 2222 3716
rect 2158 2930 2164 3712
rect 2216 2930 2222 3712
rect 1849 2922 1895 2926
rect 2007 2922 2053 2928
rect 2158 2926 2222 2930
rect 2316 3714 2380 3718
rect 2481 3716 2527 3722
rect 2639 3718 2685 3722
rect 2316 2932 2322 3714
rect 2374 2932 2380 3714
rect 2316 2928 2380 2932
rect 2474 3712 2538 3716
rect 2474 2930 2480 3712
rect 2532 2930 2538 3712
rect 2165 2922 2211 2926
rect 2323 2922 2369 2928
rect 2474 2926 2538 2930
rect 2632 3714 2696 3718
rect 2797 3716 2843 3722
rect 2955 3718 3001 3722
rect 2632 2932 2638 3714
rect 2690 2932 2696 3714
rect 2632 2928 2696 2932
rect 2790 3712 2854 3716
rect 2790 2930 2796 3712
rect 2848 2930 2854 3712
rect 2481 2922 2527 2926
rect 2639 2922 2685 2928
rect 2790 2926 2854 2930
rect 2948 3714 3012 3718
rect 3113 3716 3159 3722
rect 3271 3718 3317 3722
rect 2948 2932 2954 3714
rect 3006 2932 3012 3714
rect 2948 2928 3012 2932
rect 3106 3712 3170 3716
rect 3106 2930 3112 3712
rect 3164 2930 3170 3712
rect 2797 2922 2843 2926
rect 2955 2922 3001 2928
rect 3106 2926 3170 2930
rect 3264 3714 3328 3718
rect 3429 3716 3475 3722
rect 3587 3718 3633 3722
rect 3264 2932 3270 3714
rect 3322 2932 3328 3714
rect 3264 2928 3328 2932
rect 3422 3712 3486 3716
rect 3422 2930 3428 3712
rect 3480 2930 3486 3712
rect 3113 2922 3159 2926
rect 3271 2922 3317 2928
rect 3422 2926 3486 2930
rect 3580 3714 3644 3718
rect 3745 3716 3791 3722
rect 3903 3718 3949 3722
rect 3580 2932 3586 3714
rect 3638 2932 3644 3714
rect 3580 2928 3644 2932
rect 3738 3712 3802 3716
rect 3738 2930 3744 3712
rect 3796 2930 3802 3712
rect 3429 2922 3475 2926
rect 3587 2922 3633 2928
rect 3738 2926 3802 2930
rect 3896 3714 3960 3718
rect 4061 3716 4107 3722
rect 4219 3718 4265 3722
rect 3896 2932 3902 3714
rect 3954 2932 3960 3714
rect 3896 2928 3960 2932
rect 4054 3712 4118 3716
rect 4054 2930 4060 3712
rect 4112 2930 4118 3712
rect 3745 2922 3791 2926
rect 3903 2922 3949 2928
rect 4054 2926 4118 2930
rect 4212 3714 4276 3718
rect 4377 3716 4423 3722
rect 4535 3718 4581 3722
rect 4212 2932 4218 3714
rect 4270 2932 4276 3714
rect 4212 2928 4276 2932
rect 4370 3712 4434 3716
rect 4370 2930 4376 3712
rect 4428 2930 4434 3712
rect 4061 2922 4107 2926
rect 4219 2922 4265 2928
rect 4370 2926 4434 2930
rect 4528 3714 4592 3718
rect 4693 3716 4739 3722
rect 4851 3718 4897 3722
rect 4528 2932 4534 3714
rect 4586 2932 4592 3714
rect 4528 2928 4592 2932
rect 4686 3712 4750 3716
rect 4686 2930 4692 3712
rect 4744 2930 4750 3712
rect 4377 2922 4423 2926
rect 4535 2922 4581 2928
rect 4686 2926 4750 2930
rect 4844 3714 4908 3718
rect 5009 3716 5055 3722
rect 5167 3718 5213 3722
rect 4844 2932 4850 3714
rect 4902 2932 4908 3714
rect 4844 2928 4908 2932
rect 5002 3712 5066 3716
rect 5002 2930 5008 3712
rect 5060 2930 5066 3712
rect 4693 2922 4739 2926
rect 4851 2922 4897 2928
rect 5002 2926 5066 2930
rect 5160 3714 5224 3718
rect 5325 3716 5371 3722
rect 5483 3718 5529 3722
rect 5160 2932 5166 3714
rect 5218 2932 5224 3714
rect 5160 2928 5224 2932
rect 5318 3712 5382 3716
rect 5318 2930 5324 3712
rect 5376 2930 5382 3712
rect 5009 2922 5055 2926
rect 5167 2922 5213 2928
rect 5318 2926 5382 2930
rect 5476 3714 5540 3718
rect 5641 3716 5687 3722
rect 5799 3718 5845 3722
rect 5476 2932 5482 3714
rect 5534 2932 5540 3714
rect 5476 2928 5540 2932
rect 5634 3712 5698 3716
rect 5634 2930 5640 3712
rect 5692 2930 5698 3712
rect 5325 2922 5371 2926
rect 5483 2922 5529 2928
rect 5634 2926 5698 2930
rect 5792 3714 5856 3718
rect 5957 3716 6003 3722
rect 6115 3718 6161 3722
rect 5792 2932 5798 3714
rect 5850 2932 5856 3714
rect 5792 2928 5856 2932
rect 5950 3712 6014 3716
rect 5950 2930 5956 3712
rect 6008 2930 6014 3712
rect 5641 2922 5687 2926
rect 5799 2922 5845 2928
rect 5950 2926 6014 2930
rect 6108 3714 6172 3718
rect 6273 3716 6319 3722
rect 6431 3718 6477 3722
rect 6108 2932 6114 3714
rect 6166 2932 6172 3714
rect 6108 2928 6172 2932
rect 6266 3712 6330 3716
rect 6266 2930 6272 3712
rect 6324 2930 6330 3712
rect 5957 2922 6003 2926
rect 6115 2922 6161 2928
rect 6266 2926 6330 2930
rect 6424 3714 6488 3718
rect 6589 3716 6635 3722
rect 6747 3718 6793 3722
rect 6424 2932 6430 3714
rect 6482 2932 6488 3714
rect 6424 2928 6488 2932
rect 6582 3712 6646 3716
rect 6582 2930 6588 3712
rect 6640 2930 6646 3712
rect 6273 2922 6319 2926
rect 6431 2922 6477 2928
rect 6582 2926 6646 2930
rect 6740 3714 6804 3718
rect 6905 3716 6951 3722
rect 7063 3718 7109 3722
rect 6740 2932 6746 3714
rect 6798 2932 6804 3714
rect 6740 2928 6804 2932
rect 6898 3712 6962 3716
rect 6898 2930 6904 3712
rect 6956 2930 6962 3712
rect 6589 2922 6635 2926
rect 6747 2922 6793 2928
rect 6898 2926 6962 2930
rect 7056 3714 7120 3718
rect 7221 3716 7267 3722
rect 7379 3718 7425 3722
rect 7056 2932 7062 3714
rect 7114 2932 7120 3714
rect 7056 2928 7120 2932
rect 7214 3712 7278 3716
rect 7214 2930 7220 3712
rect 7272 2930 7278 3712
rect 6905 2922 6951 2926
rect 7063 2922 7109 2928
rect 7214 2926 7278 2930
rect 7372 3714 7436 3718
rect 7537 3716 7583 3722
rect 7695 3718 7741 3722
rect 7372 2932 7378 3714
rect 7430 2932 7436 3714
rect 7372 2928 7436 2932
rect 7530 3712 7594 3716
rect 7530 2930 7536 3712
rect 7588 2930 7594 3712
rect 7221 2922 7267 2926
rect 7379 2922 7425 2928
rect 7530 2926 7594 2930
rect 7688 3714 7752 3718
rect 7853 3716 7899 3722
rect 8011 3718 8057 3722
rect 7688 2932 7694 3714
rect 7746 2932 7752 3714
rect 7688 2928 7752 2932
rect 7846 3712 7910 3716
rect 7846 2930 7852 3712
rect 7904 2930 7910 3712
rect 7537 2922 7583 2926
rect 7695 2922 7741 2928
rect 7846 2926 7910 2930
rect 8004 3714 8068 3718
rect 8169 3716 8215 3722
rect 8327 3718 8373 3722
rect 8004 2932 8010 3714
rect 8062 2932 8068 3714
rect 8004 2928 8068 2932
rect 8162 3712 8226 3716
rect 8162 2930 8168 3712
rect 8220 2930 8226 3712
rect 7853 2922 7899 2926
rect 8011 2922 8057 2928
rect 8162 2926 8226 2930
rect 8320 3714 8384 3718
rect 8485 3716 8531 3722
rect 8643 3718 8689 3722
rect 8320 2932 8326 3714
rect 8378 2932 8384 3714
rect 8320 2928 8384 2932
rect 8478 3712 8542 3716
rect 8478 2930 8484 3712
rect 8536 2930 8542 3712
rect 8169 2922 8215 2926
rect 8327 2922 8373 2928
rect 8478 2926 8542 2930
rect 8636 3714 8700 3718
rect 8801 3716 8847 3722
rect 8959 3718 9005 3722
rect 8636 2932 8642 3714
rect 8694 2932 8700 3714
rect 8636 2928 8700 2932
rect 8794 3712 8858 3716
rect 8794 2930 8800 3712
rect 8852 2930 8858 3712
rect 8485 2922 8531 2926
rect 8643 2922 8689 2928
rect 8794 2926 8858 2930
rect 8952 3714 9016 3718
rect 9117 3716 9163 3722
rect 9275 3718 9321 3722
rect 8952 2932 8958 3714
rect 9010 2932 9016 3714
rect 8952 2928 9016 2932
rect 9110 3712 9174 3716
rect 9110 2930 9116 3712
rect 9168 2930 9174 3712
rect 8801 2922 8847 2926
rect 8959 2922 9005 2928
rect 9110 2926 9174 2930
rect 9268 3714 9332 3718
rect 9433 3716 9479 3722
rect 9591 3718 9637 3722
rect 9268 2932 9274 3714
rect 9326 2932 9332 3714
rect 9268 2928 9332 2932
rect 9426 3712 9490 3716
rect 9426 2930 9432 3712
rect 9484 2930 9490 3712
rect 9117 2922 9163 2926
rect 9275 2922 9321 2928
rect 9426 2926 9490 2930
rect 9584 3714 9648 3718
rect 9749 3716 9795 3722
rect 9907 3718 9953 3722
rect 9584 2932 9590 3714
rect 9642 2932 9648 3714
rect 9584 2928 9648 2932
rect 9742 3712 9806 3716
rect 9742 2930 9748 3712
rect 9800 2930 9806 3712
rect 9433 2922 9479 2926
rect 9591 2922 9637 2928
rect 9742 2926 9806 2930
rect 9900 3714 9964 3718
rect 10065 3716 10111 3722
rect 10223 3718 10269 3722
rect 9900 2932 9906 3714
rect 9958 2932 9964 3714
rect 9900 2928 9964 2932
rect 10058 3712 10122 3716
rect 10058 2930 10064 3712
rect 10116 2930 10122 3712
rect 9749 2922 9795 2926
rect 9907 2922 9953 2928
rect 10058 2926 10122 2930
rect 10216 3714 10280 3718
rect 10381 3716 10427 3722
rect 10539 3718 10585 3722
rect 10216 2932 10222 3714
rect 10274 2932 10280 3714
rect 10216 2928 10280 2932
rect 10374 3712 10438 3716
rect 10374 2930 10380 3712
rect 10432 2930 10438 3712
rect 10065 2922 10111 2926
rect 10223 2922 10269 2928
rect 10374 2926 10438 2930
rect 10532 3714 10596 3718
rect 10697 3716 10743 3722
rect 10855 3718 10901 3722
rect 10532 2932 10538 3714
rect 10590 2932 10596 3714
rect 10532 2928 10596 2932
rect 10690 3712 10754 3716
rect 10690 2930 10696 3712
rect 10748 2930 10754 3712
rect 10381 2922 10427 2926
rect 10539 2922 10585 2928
rect 10690 2926 10754 2930
rect 10848 3714 10912 3718
rect 11013 3716 11059 3722
rect 11171 3718 11217 3722
rect 10848 2932 10854 3714
rect 10906 2932 10912 3714
rect 10848 2928 10912 2932
rect 11006 3712 11070 3716
rect 11006 2930 11012 3712
rect 11064 2930 11070 3712
rect 10697 2922 10743 2926
rect 10855 2922 10901 2928
rect 11006 2926 11070 2930
rect 11164 3714 11228 3718
rect 11329 3716 11375 3722
rect 11487 3718 11533 3722
rect 11164 2932 11170 3714
rect 11222 2932 11228 3714
rect 11164 2928 11228 2932
rect 11322 3712 11386 3716
rect 11322 2930 11328 3712
rect 11380 2930 11386 3712
rect 11013 2922 11059 2926
rect 11171 2922 11217 2928
rect 11322 2926 11386 2930
rect 11480 3714 11544 3718
rect 11645 3716 11691 3722
rect 11803 3718 11849 3722
rect 11480 2932 11486 3714
rect 11538 2932 11544 3714
rect 11480 2928 11544 2932
rect 11638 3712 11702 3716
rect 11638 2930 11644 3712
rect 11696 2930 11702 3712
rect 11329 2922 11375 2926
rect 11487 2922 11533 2928
rect 11638 2926 11702 2930
rect 11796 3714 11860 3718
rect 11961 3716 12007 3722
rect 12119 3718 12165 3722
rect 11796 2932 11802 3714
rect 11854 2932 11860 3714
rect 11796 2928 11860 2932
rect 11954 3712 12018 3716
rect 11954 2930 11960 3712
rect 12012 2930 12018 3712
rect 11645 2922 11691 2926
rect 11803 2922 11849 2928
rect 11954 2926 12018 2930
rect 12112 3714 12176 3718
rect 12277 3716 12323 3722
rect 12435 3718 12481 3722
rect 12112 2932 12118 3714
rect 12170 2932 12176 3714
rect 12112 2928 12176 2932
rect 12270 3712 12334 3716
rect 12270 2930 12276 3712
rect 12328 2930 12334 3712
rect 11961 2922 12007 2926
rect 12119 2922 12165 2928
rect 12270 2926 12334 2930
rect 12428 3714 12492 3718
rect 12593 3716 12639 3722
rect 12745 3718 12791 3722
rect 12428 2932 12434 3714
rect 12486 2932 12492 3714
rect 12428 2928 12492 2932
rect 12586 3712 12650 3716
rect 12586 2930 12592 3712
rect 12644 2930 12650 3712
rect 12277 2922 12323 2926
rect 12435 2922 12481 2928
rect 12586 2926 12650 2930
rect 12738 3714 12802 3718
rect 12738 2932 12744 3714
rect 12796 2932 12802 3714
rect 12738 2928 12802 2932
rect 12593 2922 12639 2926
rect 12745 2922 12791 2928
rect 12830 2890 12864 3754
rect 42 2844 12864 2890
rect 12892 2894 12904 4808
rect 12938 2894 12950 4828
rect 12892 2854 12950 2894
rect 42 2712 76 2844
rect -124 2112 76 2712
rect 42 1980 76 2112
rect 104 2804 168 2808
rect 269 2806 315 2812
rect 427 2808 473 2812
rect 104 2022 110 2804
rect 162 2022 168 2804
rect 104 2018 168 2022
rect 262 2802 326 2806
rect 262 2020 268 2802
rect 320 2020 326 2802
rect 262 2016 326 2020
rect 420 2804 484 2808
rect 585 2806 631 2812
rect 743 2808 789 2812
rect 420 2022 426 2804
rect 478 2022 484 2804
rect 420 2018 484 2022
rect 578 2802 642 2806
rect 578 2020 584 2802
rect 636 2020 642 2802
rect 269 2012 315 2016
rect 427 2012 473 2018
rect 578 2016 642 2020
rect 736 2804 800 2808
rect 901 2806 947 2812
rect 1059 2808 1105 2812
rect 736 2022 742 2804
rect 794 2022 800 2804
rect 736 2018 800 2022
rect 894 2802 958 2806
rect 894 2020 900 2802
rect 952 2020 958 2802
rect 585 2012 631 2016
rect 743 2012 789 2018
rect 894 2016 958 2020
rect 1052 2804 1116 2808
rect 1217 2806 1263 2812
rect 1375 2808 1421 2812
rect 1052 2022 1058 2804
rect 1110 2022 1116 2804
rect 1052 2018 1116 2022
rect 1210 2802 1274 2806
rect 1210 2020 1216 2802
rect 1268 2020 1274 2802
rect 901 2012 947 2016
rect 1059 2012 1105 2018
rect 1210 2016 1274 2020
rect 1368 2804 1432 2808
rect 1533 2806 1579 2812
rect 1691 2808 1737 2812
rect 1368 2022 1374 2804
rect 1426 2022 1432 2804
rect 1368 2018 1432 2022
rect 1526 2802 1590 2806
rect 1526 2020 1532 2802
rect 1584 2020 1590 2802
rect 1217 2012 1263 2016
rect 1375 2012 1421 2018
rect 1526 2016 1590 2020
rect 1684 2804 1748 2808
rect 1849 2806 1895 2812
rect 2007 2808 2053 2812
rect 1684 2022 1690 2804
rect 1742 2022 1748 2804
rect 1684 2018 1748 2022
rect 1842 2802 1906 2806
rect 1842 2020 1848 2802
rect 1900 2020 1906 2802
rect 1533 2012 1579 2016
rect 1691 2012 1737 2018
rect 1842 2016 1906 2020
rect 2000 2804 2064 2808
rect 2165 2806 2211 2812
rect 2323 2808 2369 2812
rect 2000 2022 2006 2804
rect 2058 2022 2064 2804
rect 2000 2018 2064 2022
rect 2158 2802 2222 2806
rect 2158 2020 2164 2802
rect 2216 2020 2222 2802
rect 1849 2012 1895 2016
rect 2007 2012 2053 2018
rect 2158 2016 2222 2020
rect 2316 2804 2380 2808
rect 2481 2806 2527 2812
rect 2639 2808 2685 2812
rect 2316 2022 2322 2804
rect 2374 2022 2380 2804
rect 2316 2018 2380 2022
rect 2474 2802 2538 2806
rect 2474 2020 2480 2802
rect 2532 2020 2538 2802
rect 2165 2012 2211 2016
rect 2323 2012 2369 2018
rect 2474 2016 2538 2020
rect 2632 2804 2696 2808
rect 2797 2806 2843 2812
rect 2955 2808 3001 2812
rect 2632 2022 2638 2804
rect 2690 2022 2696 2804
rect 2632 2018 2696 2022
rect 2790 2802 2854 2806
rect 2790 2020 2796 2802
rect 2848 2020 2854 2802
rect 2481 2012 2527 2016
rect 2639 2012 2685 2018
rect 2790 2016 2854 2020
rect 2948 2804 3012 2808
rect 3113 2806 3159 2812
rect 3271 2808 3317 2812
rect 2948 2022 2954 2804
rect 3006 2022 3012 2804
rect 2948 2018 3012 2022
rect 3106 2802 3170 2806
rect 3106 2020 3112 2802
rect 3164 2020 3170 2802
rect 2797 2012 2843 2016
rect 2955 2012 3001 2018
rect 3106 2016 3170 2020
rect 3264 2804 3328 2808
rect 3429 2806 3475 2812
rect 3587 2808 3633 2812
rect 3264 2022 3270 2804
rect 3322 2022 3328 2804
rect 3264 2018 3328 2022
rect 3422 2802 3486 2806
rect 3422 2020 3428 2802
rect 3480 2020 3486 2802
rect 3113 2012 3159 2016
rect 3271 2012 3317 2018
rect 3422 2016 3486 2020
rect 3580 2804 3644 2808
rect 3745 2806 3791 2812
rect 3903 2808 3949 2812
rect 3580 2022 3586 2804
rect 3638 2022 3644 2804
rect 3580 2018 3644 2022
rect 3738 2802 3802 2806
rect 3738 2020 3744 2802
rect 3796 2020 3802 2802
rect 3429 2012 3475 2016
rect 3587 2012 3633 2018
rect 3738 2016 3802 2020
rect 3896 2804 3960 2808
rect 4061 2806 4107 2812
rect 4219 2808 4265 2812
rect 3896 2022 3902 2804
rect 3954 2022 3960 2804
rect 3896 2018 3960 2022
rect 4054 2802 4118 2806
rect 4054 2020 4060 2802
rect 4112 2020 4118 2802
rect 3745 2012 3791 2016
rect 3903 2012 3949 2018
rect 4054 2016 4118 2020
rect 4212 2804 4276 2808
rect 4377 2806 4423 2812
rect 4535 2808 4581 2812
rect 4212 2022 4218 2804
rect 4270 2022 4276 2804
rect 4212 2018 4276 2022
rect 4370 2802 4434 2806
rect 4370 2020 4376 2802
rect 4428 2020 4434 2802
rect 4061 2012 4107 2016
rect 4219 2012 4265 2018
rect 4370 2016 4434 2020
rect 4528 2804 4592 2808
rect 4693 2806 4739 2812
rect 4851 2808 4897 2812
rect 4528 2022 4534 2804
rect 4586 2022 4592 2804
rect 4528 2018 4592 2022
rect 4686 2802 4750 2806
rect 4686 2020 4692 2802
rect 4744 2020 4750 2802
rect 4377 2012 4423 2016
rect 4535 2012 4581 2018
rect 4686 2016 4750 2020
rect 4844 2804 4908 2808
rect 5009 2806 5055 2812
rect 5167 2808 5213 2812
rect 4844 2022 4850 2804
rect 4902 2022 4908 2804
rect 4844 2018 4908 2022
rect 5002 2802 5066 2806
rect 5002 2020 5008 2802
rect 5060 2020 5066 2802
rect 4693 2012 4739 2016
rect 4851 2012 4897 2018
rect 5002 2016 5066 2020
rect 5160 2804 5224 2808
rect 5325 2806 5371 2812
rect 5483 2808 5529 2812
rect 5160 2022 5166 2804
rect 5218 2022 5224 2804
rect 5160 2018 5224 2022
rect 5318 2802 5382 2806
rect 5318 2020 5324 2802
rect 5376 2020 5382 2802
rect 5009 2012 5055 2016
rect 5167 2012 5213 2018
rect 5318 2016 5382 2020
rect 5476 2804 5540 2808
rect 5641 2806 5687 2812
rect 5799 2808 5845 2812
rect 5476 2022 5482 2804
rect 5534 2022 5540 2804
rect 5476 2018 5540 2022
rect 5634 2802 5698 2806
rect 5634 2020 5640 2802
rect 5692 2020 5698 2802
rect 5325 2012 5371 2016
rect 5483 2012 5529 2018
rect 5634 2016 5698 2020
rect 5792 2804 5856 2808
rect 5957 2806 6003 2812
rect 6115 2808 6161 2812
rect 5792 2022 5798 2804
rect 5850 2022 5856 2804
rect 5792 2018 5856 2022
rect 5950 2802 6014 2806
rect 5950 2020 5956 2802
rect 6008 2020 6014 2802
rect 5641 2012 5687 2016
rect 5799 2012 5845 2018
rect 5950 2016 6014 2020
rect 6108 2804 6172 2808
rect 6273 2806 6319 2812
rect 6431 2808 6477 2812
rect 6108 2022 6114 2804
rect 6166 2022 6172 2804
rect 6108 2018 6172 2022
rect 6266 2802 6330 2806
rect 6266 2020 6272 2802
rect 6324 2020 6330 2802
rect 5957 2012 6003 2016
rect 6115 2012 6161 2018
rect 6266 2016 6330 2020
rect 6424 2804 6488 2808
rect 6589 2806 6635 2812
rect 6747 2808 6793 2812
rect 6424 2022 6430 2804
rect 6482 2022 6488 2804
rect 6424 2018 6488 2022
rect 6582 2802 6646 2806
rect 6582 2020 6588 2802
rect 6640 2020 6646 2802
rect 6273 2012 6319 2016
rect 6431 2012 6477 2018
rect 6582 2016 6646 2020
rect 6740 2804 6804 2808
rect 6905 2806 6951 2812
rect 7063 2808 7109 2812
rect 6740 2022 6746 2804
rect 6798 2022 6804 2804
rect 6740 2018 6804 2022
rect 6898 2802 6962 2806
rect 6898 2020 6904 2802
rect 6956 2020 6962 2802
rect 6589 2012 6635 2016
rect 6747 2012 6793 2018
rect 6898 2016 6962 2020
rect 7056 2804 7120 2808
rect 7221 2806 7267 2812
rect 7379 2808 7425 2812
rect 7056 2022 7062 2804
rect 7114 2022 7120 2804
rect 7056 2018 7120 2022
rect 7214 2802 7278 2806
rect 7214 2020 7220 2802
rect 7272 2020 7278 2802
rect 6905 2012 6951 2016
rect 7063 2012 7109 2018
rect 7214 2016 7278 2020
rect 7372 2804 7436 2808
rect 7537 2806 7583 2812
rect 7695 2808 7741 2812
rect 7372 2022 7378 2804
rect 7430 2022 7436 2804
rect 7372 2018 7436 2022
rect 7530 2802 7594 2806
rect 7530 2020 7536 2802
rect 7588 2020 7594 2802
rect 7221 2012 7267 2016
rect 7379 2012 7425 2018
rect 7530 2016 7594 2020
rect 7688 2804 7752 2808
rect 7853 2806 7899 2812
rect 8011 2808 8057 2812
rect 7688 2022 7694 2804
rect 7746 2022 7752 2804
rect 7688 2018 7752 2022
rect 7846 2802 7910 2806
rect 7846 2020 7852 2802
rect 7904 2020 7910 2802
rect 7537 2012 7583 2016
rect 7695 2012 7741 2018
rect 7846 2016 7910 2020
rect 8004 2804 8068 2808
rect 8169 2806 8215 2812
rect 8327 2808 8373 2812
rect 8004 2022 8010 2804
rect 8062 2022 8068 2804
rect 8004 2018 8068 2022
rect 8162 2802 8226 2806
rect 8162 2020 8168 2802
rect 8220 2020 8226 2802
rect 7853 2012 7899 2016
rect 8011 2012 8057 2018
rect 8162 2016 8226 2020
rect 8320 2804 8384 2808
rect 8485 2806 8531 2812
rect 8643 2808 8689 2812
rect 8320 2022 8326 2804
rect 8378 2022 8384 2804
rect 8320 2018 8384 2022
rect 8478 2802 8542 2806
rect 8478 2020 8484 2802
rect 8536 2020 8542 2802
rect 8169 2012 8215 2016
rect 8327 2012 8373 2018
rect 8478 2016 8542 2020
rect 8636 2804 8700 2808
rect 8801 2806 8847 2812
rect 8959 2808 9005 2812
rect 8636 2022 8642 2804
rect 8694 2022 8700 2804
rect 8636 2018 8700 2022
rect 8794 2802 8858 2806
rect 8794 2020 8800 2802
rect 8852 2020 8858 2802
rect 8485 2012 8531 2016
rect 8643 2012 8689 2018
rect 8794 2016 8858 2020
rect 8952 2804 9016 2808
rect 9117 2806 9163 2812
rect 9275 2808 9321 2812
rect 8952 2022 8958 2804
rect 9010 2022 9016 2804
rect 8952 2018 9016 2022
rect 9110 2802 9174 2806
rect 9110 2020 9116 2802
rect 9168 2020 9174 2802
rect 8801 2012 8847 2016
rect 8959 2012 9005 2018
rect 9110 2016 9174 2020
rect 9268 2804 9332 2808
rect 9433 2806 9479 2812
rect 9591 2808 9637 2812
rect 9268 2022 9274 2804
rect 9326 2022 9332 2804
rect 9268 2018 9332 2022
rect 9426 2802 9490 2806
rect 9426 2020 9432 2802
rect 9484 2020 9490 2802
rect 9117 2012 9163 2016
rect 9275 2012 9321 2018
rect 9426 2016 9490 2020
rect 9584 2804 9648 2808
rect 9749 2806 9795 2812
rect 9907 2808 9953 2812
rect 9584 2022 9590 2804
rect 9642 2022 9648 2804
rect 9584 2018 9648 2022
rect 9742 2802 9806 2806
rect 9742 2020 9748 2802
rect 9800 2020 9806 2802
rect 9433 2012 9479 2016
rect 9591 2012 9637 2018
rect 9742 2016 9806 2020
rect 9900 2804 9964 2808
rect 10065 2806 10111 2812
rect 10223 2808 10269 2812
rect 9900 2022 9906 2804
rect 9958 2022 9964 2804
rect 9900 2018 9964 2022
rect 10058 2802 10122 2806
rect 10058 2020 10064 2802
rect 10116 2020 10122 2802
rect 9749 2012 9795 2016
rect 9907 2012 9953 2018
rect 10058 2016 10122 2020
rect 10216 2804 10280 2808
rect 10381 2806 10427 2812
rect 10539 2808 10585 2812
rect 10216 2022 10222 2804
rect 10274 2022 10280 2804
rect 10216 2018 10280 2022
rect 10374 2802 10438 2806
rect 10374 2020 10380 2802
rect 10432 2020 10438 2802
rect 10065 2012 10111 2016
rect 10223 2012 10269 2018
rect 10374 2016 10438 2020
rect 10532 2804 10596 2808
rect 10697 2806 10743 2812
rect 10855 2808 10901 2812
rect 10532 2022 10538 2804
rect 10590 2022 10596 2804
rect 10532 2018 10596 2022
rect 10690 2802 10754 2806
rect 10690 2020 10696 2802
rect 10748 2020 10754 2802
rect 10381 2012 10427 2016
rect 10539 2012 10585 2018
rect 10690 2016 10754 2020
rect 10848 2804 10912 2808
rect 11013 2806 11059 2812
rect 11171 2808 11217 2812
rect 10848 2022 10854 2804
rect 10906 2022 10912 2804
rect 10848 2018 10912 2022
rect 11006 2802 11070 2806
rect 11006 2020 11012 2802
rect 11064 2020 11070 2802
rect 10697 2012 10743 2016
rect 10855 2012 10901 2018
rect 11006 2016 11070 2020
rect 11164 2804 11228 2808
rect 11329 2806 11375 2812
rect 11487 2808 11533 2812
rect 11164 2022 11170 2804
rect 11222 2022 11228 2804
rect 11164 2018 11228 2022
rect 11322 2802 11386 2806
rect 11322 2020 11328 2802
rect 11380 2020 11386 2802
rect 11013 2012 11059 2016
rect 11171 2012 11217 2018
rect 11322 2016 11386 2020
rect 11480 2804 11544 2808
rect 11645 2806 11691 2812
rect 11803 2808 11849 2812
rect 11480 2022 11486 2804
rect 11538 2022 11544 2804
rect 11480 2018 11544 2022
rect 11638 2802 11702 2806
rect 11638 2020 11644 2802
rect 11696 2020 11702 2802
rect 11329 2012 11375 2016
rect 11487 2012 11533 2018
rect 11638 2016 11702 2020
rect 11796 2804 11860 2808
rect 11961 2806 12007 2812
rect 12119 2808 12165 2812
rect 11796 2022 11802 2804
rect 11854 2022 11860 2804
rect 11796 2018 11860 2022
rect 11954 2802 12018 2806
rect 11954 2020 11960 2802
rect 12012 2020 12018 2802
rect 11645 2012 11691 2016
rect 11803 2012 11849 2018
rect 11954 2016 12018 2020
rect 12112 2804 12176 2808
rect 12277 2806 12323 2812
rect 12435 2808 12481 2812
rect 12112 2022 12118 2804
rect 12170 2022 12176 2804
rect 12112 2018 12176 2022
rect 12270 2802 12334 2806
rect 12270 2020 12276 2802
rect 12328 2020 12334 2802
rect 11961 2012 12007 2016
rect 12119 2012 12165 2018
rect 12270 2016 12334 2020
rect 12428 2804 12492 2808
rect 12593 2806 12639 2812
rect 12745 2808 12791 2812
rect 12428 2022 12434 2804
rect 12486 2022 12492 2804
rect 12428 2018 12492 2022
rect 12586 2802 12650 2806
rect 12586 2020 12592 2802
rect 12644 2020 12650 2802
rect 12277 2012 12323 2016
rect 12435 2012 12481 2018
rect 12586 2016 12650 2020
rect 12738 2804 12802 2808
rect 12738 2022 12744 2804
rect 12796 2022 12802 2804
rect 12738 2018 12802 2022
rect 12830 2712 12864 2844
rect 12830 2112 13030 2712
rect 12593 2012 12639 2016
rect 12745 2012 12791 2018
rect 12830 1980 12864 2112
rect -44 1932 14 1972
rect -44 -6 -32 1932
rect 2 16 14 1932
rect 42 1934 12864 1980
rect 42 1070 76 1934
rect 104 1894 168 1898
rect 269 1896 315 1902
rect 427 1898 473 1902
rect 104 1112 110 1894
rect 162 1112 168 1894
rect 104 1108 168 1112
rect 262 1892 326 1896
rect 262 1110 268 1892
rect 320 1110 326 1892
rect 262 1106 326 1110
rect 420 1894 484 1898
rect 585 1896 631 1902
rect 743 1898 789 1902
rect 420 1112 426 1894
rect 478 1112 484 1894
rect 420 1108 484 1112
rect 578 1892 642 1896
rect 578 1110 584 1892
rect 636 1110 642 1892
rect 269 1102 315 1106
rect 427 1102 473 1108
rect 578 1106 642 1110
rect 736 1894 800 1898
rect 901 1896 947 1902
rect 1059 1898 1105 1902
rect 736 1112 742 1894
rect 794 1112 800 1894
rect 736 1108 800 1112
rect 894 1892 958 1896
rect 894 1110 900 1892
rect 952 1110 958 1892
rect 585 1102 631 1106
rect 743 1102 789 1108
rect 894 1106 958 1110
rect 1052 1894 1116 1898
rect 1217 1896 1263 1902
rect 1375 1898 1421 1902
rect 1052 1112 1058 1894
rect 1110 1112 1116 1894
rect 1052 1108 1116 1112
rect 1210 1892 1274 1896
rect 1210 1110 1216 1892
rect 1268 1110 1274 1892
rect 901 1102 947 1106
rect 1059 1102 1105 1108
rect 1210 1106 1274 1110
rect 1368 1894 1432 1898
rect 1533 1896 1579 1902
rect 1691 1898 1737 1902
rect 1368 1112 1374 1894
rect 1426 1112 1432 1894
rect 1368 1108 1432 1112
rect 1526 1892 1590 1896
rect 1526 1110 1532 1892
rect 1584 1110 1590 1892
rect 1217 1102 1263 1106
rect 1375 1102 1421 1108
rect 1526 1106 1590 1110
rect 1684 1894 1748 1898
rect 1849 1896 1895 1902
rect 2007 1898 2053 1902
rect 1684 1112 1690 1894
rect 1742 1112 1748 1894
rect 1684 1108 1748 1112
rect 1842 1892 1906 1896
rect 1842 1110 1848 1892
rect 1900 1110 1906 1892
rect 1533 1102 1579 1106
rect 1691 1102 1737 1108
rect 1842 1106 1906 1110
rect 2000 1894 2064 1898
rect 2165 1896 2211 1902
rect 2323 1898 2369 1902
rect 2000 1112 2006 1894
rect 2058 1112 2064 1894
rect 2000 1108 2064 1112
rect 2158 1892 2222 1896
rect 2158 1110 2164 1892
rect 2216 1110 2222 1892
rect 1849 1102 1895 1106
rect 2007 1102 2053 1108
rect 2158 1106 2222 1110
rect 2316 1894 2380 1898
rect 2481 1896 2527 1902
rect 2639 1898 2685 1902
rect 2316 1112 2322 1894
rect 2374 1112 2380 1894
rect 2316 1108 2380 1112
rect 2474 1892 2538 1896
rect 2474 1110 2480 1892
rect 2532 1110 2538 1892
rect 2165 1102 2211 1106
rect 2323 1102 2369 1108
rect 2474 1106 2538 1110
rect 2632 1894 2696 1898
rect 2797 1896 2843 1902
rect 2955 1898 3001 1902
rect 2632 1112 2638 1894
rect 2690 1112 2696 1894
rect 2632 1108 2696 1112
rect 2790 1892 2854 1896
rect 2790 1110 2796 1892
rect 2848 1110 2854 1892
rect 2481 1102 2527 1106
rect 2639 1102 2685 1108
rect 2790 1106 2854 1110
rect 2948 1894 3012 1898
rect 3113 1896 3159 1902
rect 3271 1898 3317 1902
rect 2948 1112 2954 1894
rect 3006 1112 3012 1894
rect 2948 1108 3012 1112
rect 3106 1892 3170 1896
rect 3106 1110 3112 1892
rect 3164 1110 3170 1892
rect 2797 1102 2843 1106
rect 2955 1102 3001 1108
rect 3106 1106 3170 1110
rect 3264 1894 3328 1898
rect 3429 1896 3475 1902
rect 3587 1898 3633 1902
rect 3264 1112 3270 1894
rect 3322 1112 3328 1894
rect 3264 1108 3328 1112
rect 3422 1892 3486 1896
rect 3422 1110 3428 1892
rect 3480 1110 3486 1892
rect 3113 1102 3159 1106
rect 3271 1102 3317 1108
rect 3422 1106 3486 1110
rect 3580 1894 3644 1898
rect 3745 1896 3791 1902
rect 3903 1898 3949 1902
rect 3580 1112 3586 1894
rect 3638 1112 3644 1894
rect 3580 1108 3644 1112
rect 3738 1892 3802 1896
rect 3738 1110 3744 1892
rect 3796 1110 3802 1892
rect 3429 1102 3475 1106
rect 3587 1102 3633 1108
rect 3738 1106 3802 1110
rect 3896 1894 3960 1898
rect 4061 1896 4107 1902
rect 4219 1898 4265 1902
rect 3896 1112 3902 1894
rect 3954 1112 3960 1894
rect 3896 1108 3960 1112
rect 4054 1892 4118 1896
rect 4054 1110 4060 1892
rect 4112 1110 4118 1892
rect 3745 1102 3791 1106
rect 3903 1102 3949 1108
rect 4054 1106 4118 1110
rect 4212 1894 4276 1898
rect 4377 1896 4423 1902
rect 4535 1898 4581 1902
rect 4212 1112 4218 1894
rect 4270 1112 4276 1894
rect 4212 1108 4276 1112
rect 4370 1892 4434 1896
rect 4370 1110 4376 1892
rect 4428 1110 4434 1892
rect 4061 1102 4107 1106
rect 4219 1102 4265 1108
rect 4370 1106 4434 1110
rect 4528 1894 4592 1898
rect 4693 1896 4739 1902
rect 4851 1898 4897 1902
rect 4528 1112 4534 1894
rect 4586 1112 4592 1894
rect 4528 1108 4592 1112
rect 4686 1892 4750 1896
rect 4686 1110 4692 1892
rect 4744 1110 4750 1892
rect 4377 1102 4423 1106
rect 4535 1102 4581 1108
rect 4686 1106 4750 1110
rect 4844 1894 4908 1898
rect 5009 1896 5055 1902
rect 5167 1898 5213 1902
rect 4844 1112 4850 1894
rect 4902 1112 4908 1894
rect 4844 1108 4908 1112
rect 5002 1892 5066 1896
rect 5002 1110 5008 1892
rect 5060 1110 5066 1892
rect 4693 1102 4739 1106
rect 4851 1102 4897 1108
rect 5002 1106 5066 1110
rect 5160 1894 5224 1898
rect 5325 1896 5371 1902
rect 5483 1898 5529 1902
rect 5160 1112 5166 1894
rect 5218 1112 5224 1894
rect 5160 1108 5224 1112
rect 5318 1892 5382 1896
rect 5318 1110 5324 1892
rect 5376 1110 5382 1892
rect 5009 1102 5055 1106
rect 5167 1102 5213 1108
rect 5318 1106 5382 1110
rect 5476 1894 5540 1898
rect 5641 1896 5687 1902
rect 5799 1898 5845 1902
rect 5476 1112 5482 1894
rect 5534 1112 5540 1894
rect 5476 1108 5540 1112
rect 5634 1892 5698 1896
rect 5634 1110 5640 1892
rect 5692 1110 5698 1892
rect 5325 1102 5371 1106
rect 5483 1102 5529 1108
rect 5634 1106 5698 1110
rect 5792 1894 5856 1898
rect 5957 1896 6003 1902
rect 6115 1898 6161 1902
rect 5792 1112 5798 1894
rect 5850 1112 5856 1894
rect 5792 1108 5856 1112
rect 5950 1892 6014 1896
rect 5950 1110 5956 1892
rect 6008 1110 6014 1892
rect 5641 1102 5687 1106
rect 5799 1102 5845 1108
rect 5950 1106 6014 1110
rect 6108 1894 6172 1898
rect 6273 1896 6319 1902
rect 6431 1898 6477 1902
rect 6108 1112 6114 1894
rect 6166 1112 6172 1894
rect 6108 1108 6172 1112
rect 6266 1892 6330 1896
rect 6266 1110 6272 1892
rect 6324 1110 6330 1892
rect 5957 1102 6003 1106
rect 6115 1102 6161 1108
rect 6266 1106 6330 1110
rect 6424 1894 6488 1898
rect 6589 1896 6635 1902
rect 6747 1898 6793 1902
rect 6424 1112 6430 1894
rect 6482 1112 6488 1894
rect 6424 1108 6488 1112
rect 6582 1892 6646 1896
rect 6582 1110 6588 1892
rect 6640 1110 6646 1892
rect 6273 1102 6319 1106
rect 6431 1102 6477 1108
rect 6582 1106 6646 1110
rect 6740 1894 6804 1898
rect 6905 1896 6951 1902
rect 7063 1898 7109 1902
rect 6740 1112 6746 1894
rect 6798 1112 6804 1894
rect 6740 1108 6804 1112
rect 6898 1892 6962 1896
rect 6898 1110 6904 1892
rect 6956 1110 6962 1892
rect 6589 1102 6635 1106
rect 6747 1102 6793 1108
rect 6898 1106 6962 1110
rect 7056 1894 7120 1898
rect 7221 1896 7267 1902
rect 7379 1898 7425 1902
rect 7056 1112 7062 1894
rect 7114 1112 7120 1894
rect 7056 1108 7120 1112
rect 7214 1892 7278 1896
rect 7214 1110 7220 1892
rect 7272 1110 7278 1892
rect 6905 1102 6951 1106
rect 7063 1102 7109 1108
rect 7214 1106 7278 1110
rect 7372 1894 7436 1898
rect 7537 1896 7583 1902
rect 7695 1898 7741 1902
rect 7372 1112 7378 1894
rect 7430 1112 7436 1894
rect 7372 1108 7436 1112
rect 7530 1892 7594 1896
rect 7530 1110 7536 1892
rect 7588 1110 7594 1892
rect 7221 1102 7267 1106
rect 7379 1102 7425 1108
rect 7530 1106 7594 1110
rect 7688 1894 7752 1898
rect 7853 1896 7899 1902
rect 8011 1898 8057 1902
rect 7688 1112 7694 1894
rect 7746 1112 7752 1894
rect 7688 1108 7752 1112
rect 7846 1892 7910 1896
rect 7846 1110 7852 1892
rect 7904 1110 7910 1892
rect 7537 1102 7583 1106
rect 7695 1102 7741 1108
rect 7846 1106 7910 1110
rect 8004 1894 8068 1898
rect 8169 1896 8215 1902
rect 8327 1898 8373 1902
rect 8004 1112 8010 1894
rect 8062 1112 8068 1894
rect 8004 1108 8068 1112
rect 8162 1892 8226 1896
rect 8162 1110 8168 1892
rect 8220 1110 8226 1892
rect 7853 1102 7899 1106
rect 8011 1102 8057 1108
rect 8162 1106 8226 1110
rect 8320 1894 8384 1898
rect 8485 1896 8531 1902
rect 8643 1898 8689 1902
rect 8320 1112 8326 1894
rect 8378 1112 8384 1894
rect 8320 1108 8384 1112
rect 8478 1892 8542 1896
rect 8478 1110 8484 1892
rect 8536 1110 8542 1892
rect 8169 1102 8215 1106
rect 8327 1102 8373 1108
rect 8478 1106 8542 1110
rect 8636 1894 8700 1898
rect 8801 1896 8847 1902
rect 8959 1898 9005 1902
rect 8636 1112 8642 1894
rect 8694 1112 8700 1894
rect 8636 1108 8700 1112
rect 8794 1892 8858 1896
rect 8794 1110 8800 1892
rect 8852 1110 8858 1892
rect 8485 1102 8531 1106
rect 8643 1102 8689 1108
rect 8794 1106 8858 1110
rect 8952 1894 9016 1898
rect 9117 1896 9163 1902
rect 9275 1898 9321 1902
rect 8952 1112 8958 1894
rect 9010 1112 9016 1894
rect 8952 1108 9016 1112
rect 9110 1892 9174 1896
rect 9110 1110 9116 1892
rect 9168 1110 9174 1892
rect 8801 1102 8847 1106
rect 8959 1102 9005 1108
rect 9110 1106 9174 1110
rect 9268 1894 9332 1898
rect 9433 1896 9479 1902
rect 9591 1898 9637 1902
rect 9268 1112 9274 1894
rect 9326 1112 9332 1894
rect 9268 1108 9332 1112
rect 9426 1892 9490 1896
rect 9426 1110 9432 1892
rect 9484 1110 9490 1892
rect 9117 1102 9163 1106
rect 9275 1102 9321 1108
rect 9426 1106 9490 1110
rect 9584 1894 9648 1898
rect 9749 1896 9795 1902
rect 9907 1898 9953 1902
rect 9584 1112 9590 1894
rect 9642 1112 9648 1894
rect 9584 1108 9648 1112
rect 9742 1892 9806 1896
rect 9742 1110 9748 1892
rect 9800 1110 9806 1892
rect 9433 1102 9479 1106
rect 9591 1102 9637 1108
rect 9742 1106 9806 1110
rect 9900 1894 9964 1898
rect 10065 1896 10111 1902
rect 10223 1898 10269 1902
rect 9900 1112 9906 1894
rect 9958 1112 9964 1894
rect 9900 1108 9964 1112
rect 10058 1892 10122 1896
rect 10058 1110 10064 1892
rect 10116 1110 10122 1892
rect 9749 1102 9795 1106
rect 9907 1102 9953 1108
rect 10058 1106 10122 1110
rect 10216 1894 10280 1898
rect 10381 1896 10427 1902
rect 10539 1898 10585 1902
rect 10216 1112 10222 1894
rect 10274 1112 10280 1894
rect 10216 1108 10280 1112
rect 10374 1892 10438 1896
rect 10374 1110 10380 1892
rect 10432 1110 10438 1892
rect 10065 1102 10111 1106
rect 10223 1102 10269 1108
rect 10374 1106 10438 1110
rect 10532 1894 10596 1898
rect 10697 1896 10743 1902
rect 10855 1898 10901 1902
rect 10532 1112 10538 1894
rect 10590 1112 10596 1894
rect 10532 1108 10596 1112
rect 10690 1892 10754 1896
rect 10690 1110 10696 1892
rect 10748 1110 10754 1892
rect 10381 1102 10427 1106
rect 10539 1102 10585 1108
rect 10690 1106 10754 1110
rect 10848 1894 10912 1898
rect 11013 1896 11059 1902
rect 11171 1898 11217 1902
rect 10848 1112 10854 1894
rect 10906 1112 10912 1894
rect 10848 1108 10912 1112
rect 11006 1892 11070 1896
rect 11006 1110 11012 1892
rect 11064 1110 11070 1892
rect 10697 1102 10743 1106
rect 10855 1102 10901 1108
rect 11006 1106 11070 1110
rect 11164 1894 11228 1898
rect 11329 1896 11375 1902
rect 11487 1898 11533 1902
rect 11164 1112 11170 1894
rect 11222 1112 11228 1894
rect 11164 1108 11228 1112
rect 11322 1892 11386 1896
rect 11322 1110 11328 1892
rect 11380 1110 11386 1892
rect 11013 1102 11059 1106
rect 11171 1102 11217 1108
rect 11322 1106 11386 1110
rect 11480 1894 11544 1898
rect 11645 1896 11691 1902
rect 11803 1898 11849 1902
rect 11480 1112 11486 1894
rect 11538 1112 11544 1894
rect 11480 1108 11544 1112
rect 11638 1892 11702 1896
rect 11638 1110 11644 1892
rect 11696 1110 11702 1892
rect 11329 1102 11375 1106
rect 11487 1102 11533 1108
rect 11638 1106 11702 1110
rect 11796 1894 11860 1898
rect 11961 1896 12007 1902
rect 12119 1898 12165 1902
rect 11796 1112 11802 1894
rect 11854 1112 11860 1894
rect 11796 1108 11860 1112
rect 11954 1892 12018 1896
rect 11954 1110 11960 1892
rect 12012 1110 12018 1892
rect 11645 1102 11691 1106
rect 11803 1102 11849 1108
rect 11954 1106 12018 1110
rect 12112 1894 12176 1898
rect 12277 1896 12323 1902
rect 12435 1898 12481 1902
rect 12112 1112 12118 1894
rect 12170 1112 12176 1894
rect 12112 1108 12176 1112
rect 12270 1892 12334 1896
rect 12270 1110 12276 1892
rect 12328 1110 12334 1892
rect 11961 1102 12007 1106
rect 12119 1102 12165 1108
rect 12270 1106 12334 1110
rect 12428 1894 12492 1898
rect 12593 1896 12639 1902
rect 12745 1898 12791 1902
rect 12428 1112 12434 1894
rect 12486 1112 12492 1894
rect 12428 1108 12492 1112
rect 12586 1892 12650 1896
rect 12586 1110 12592 1892
rect 12644 1110 12650 1892
rect 12277 1102 12323 1106
rect 12435 1102 12481 1108
rect 12586 1106 12650 1110
rect 12738 1894 12802 1898
rect 12738 1112 12744 1894
rect 12796 1112 12802 1894
rect 12738 1108 12802 1112
rect 12593 1102 12639 1106
rect 12745 1102 12791 1108
rect 12830 1070 12864 1934
rect 42 1024 12864 1070
rect 42 160 76 1024
rect 104 984 168 988
rect 269 986 315 992
rect 427 988 473 992
rect 104 202 110 984
rect 162 202 168 984
rect 104 198 168 202
rect 262 980 326 986
rect 262 202 268 980
rect 320 202 326 980
rect 262 196 326 202
rect 420 984 484 988
rect 585 986 631 992
rect 743 988 789 992
rect 420 202 426 984
rect 478 202 484 984
rect 420 198 484 202
rect 578 980 642 986
rect 578 202 584 980
rect 636 202 642 980
rect 269 192 315 196
rect 427 192 473 198
rect 578 196 642 202
rect 736 984 800 988
rect 901 986 947 992
rect 1059 988 1105 992
rect 736 202 742 984
rect 794 202 800 984
rect 736 198 800 202
rect 894 980 958 986
rect 894 202 900 980
rect 952 202 958 980
rect 585 192 631 196
rect 743 192 789 198
rect 894 196 958 202
rect 1052 984 1116 988
rect 1217 986 1263 992
rect 1375 988 1421 992
rect 1052 202 1058 984
rect 1110 202 1116 984
rect 1052 198 1116 202
rect 1210 980 1274 986
rect 1210 202 1216 980
rect 1268 202 1274 980
rect 901 192 947 196
rect 1059 192 1105 198
rect 1210 196 1274 202
rect 1368 984 1432 988
rect 1533 986 1579 992
rect 1691 988 1737 992
rect 1368 202 1374 984
rect 1426 202 1432 984
rect 1368 198 1432 202
rect 1526 980 1590 986
rect 1526 202 1532 980
rect 1584 202 1590 980
rect 1217 192 1263 196
rect 1375 192 1421 198
rect 1526 196 1590 202
rect 1684 984 1748 988
rect 1849 986 1895 992
rect 2007 988 2053 992
rect 1684 202 1690 984
rect 1742 202 1748 984
rect 1684 198 1748 202
rect 1842 980 1906 986
rect 1842 202 1848 980
rect 1900 202 1906 980
rect 1533 192 1579 196
rect 1691 192 1737 198
rect 1842 196 1906 202
rect 2000 984 2064 988
rect 2165 986 2211 992
rect 2323 988 2369 992
rect 2000 202 2006 984
rect 2058 202 2064 984
rect 2000 198 2064 202
rect 2158 980 2222 986
rect 2158 202 2164 980
rect 2216 202 2222 980
rect 1849 192 1895 196
rect 2007 192 2053 198
rect 2158 196 2222 202
rect 2316 984 2380 988
rect 2481 986 2527 992
rect 2639 988 2685 992
rect 2316 202 2322 984
rect 2374 202 2380 984
rect 2316 198 2380 202
rect 2474 980 2538 986
rect 2474 202 2480 980
rect 2532 202 2538 980
rect 2165 192 2211 196
rect 2323 192 2369 198
rect 2474 196 2538 202
rect 2632 984 2696 988
rect 2797 986 2843 992
rect 2955 988 3001 992
rect 2632 202 2638 984
rect 2690 202 2696 984
rect 2632 198 2696 202
rect 2790 980 2854 986
rect 2790 202 2796 980
rect 2848 202 2854 980
rect 2481 192 2527 196
rect 2639 192 2685 198
rect 2790 196 2854 202
rect 2948 984 3012 988
rect 3113 986 3159 992
rect 3271 988 3317 992
rect 2948 202 2954 984
rect 3006 202 3012 984
rect 2948 198 3012 202
rect 3106 980 3170 986
rect 3106 202 3112 980
rect 3164 202 3170 980
rect 2797 192 2843 196
rect 2955 192 3001 198
rect 3106 196 3170 202
rect 3264 984 3328 988
rect 3429 986 3475 992
rect 3587 988 3633 992
rect 3264 202 3270 984
rect 3322 202 3328 984
rect 3264 198 3328 202
rect 3422 980 3486 986
rect 3422 202 3428 980
rect 3480 202 3486 980
rect 3113 192 3159 196
rect 3271 192 3317 198
rect 3422 196 3486 202
rect 3580 984 3644 988
rect 3745 986 3791 992
rect 3903 988 3949 992
rect 3580 202 3586 984
rect 3638 202 3644 984
rect 3580 198 3644 202
rect 3738 980 3802 986
rect 3738 202 3744 980
rect 3796 202 3802 980
rect 3429 192 3475 196
rect 3587 192 3633 198
rect 3738 196 3802 202
rect 3896 984 3960 988
rect 4061 986 4107 992
rect 4219 988 4265 992
rect 3896 202 3902 984
rect 3954 202 3960 984
rect 3896 198 3960 202
rect 4054 980 4118 986
rect 4054 202 4060 980
rect 4112 202 4118 980
rect 3745 192 3791 196
rect 3903 192 3949 198
rect 4054 196 4118 202
rect 4212 984 4276 988
rect 4377 986 4423 992
rect 4535 988 4581 992
rect 4212 202 4218 984
rect 4270 202 4276 984
rect 4212 198 4276 202
rect 4370 980 4434 986
rect 4370 202 4376 980
rect 4428 202 4434 980
rect 4061 192 4107 196
rect 4219 192 4265 198
rect 4370 196 4434 202
rect 4528 984 4592 988
rect 4693 986 4739 992
rect 4851 988 4897 992
rect 4528 202 4534 984
rect 4586 202 4592 984
rect 4528 198 4592 202
rect 4686 980 4750 986
rect 4686 202 4692 980
rect 4744 202 4750 980
rect 4377 192 4423 196
rect 4535 192 4581 198
rect 4686 196 4750 202
rect 4844 984 4908 988
rect 5009 986 5055 992
rect 5167 988 5213 992
rect 4844 202 4850 984
rect 4902 202 4908 984
rect 4844 198 4908 202
rect 5002 980 5066 986
rect 5002 202 5008 980
rect 5060 202 5066 980
rect 4693 192 4739 196
rect 4851 192 4897 198
rect 5002 196 5066 202
rect 5160 984 5224 988
rect 5325 986 5371 992
rect 5483 988 5529 992
rect 5160 202 5166 984
rect 5218 202 5224 984
rect 5160 198 5224 202
rect 5318 980 5382 986
rect 5318 202 5324 980
rect 5376 202 5382 980
rect 5009 192 5055 196
rect 5167 192 5213 198
rect 5318 196 5382 202
rect 5476 984 5540 988
rect 5641 986 5687 992
rect 5799 988 5845 992
rect 5476 202 5482 984
rect 5534 202 5540 984
rect 5476 198 5540 202
rect 5634 980 5698 986
rect 5634 202 5640 980
rect 5692 202 5698 980
rect 5325 192 5371 196
rect 5483 192 5529 198
rect 5634 196 5698 202
rect 5792 984 5856 988
rect 5957 986 6003 992
rect 6115 988 6161 992
rect 5792 202 5798 984
rect 5850 202 5856 984
rect 5792 198 5856 202
rect 5950 980 6014 986
rect 5950 202 5956 980
rect 6008 202 6014 980
rect 5641 192 5687 196
rect 5799 192 5845 198
rect 5950 196 6014 202
rect 6108 984 6172 988
rect 6273 986 6319 992
rect 6431 988 6477 992
rect 6108 202 6114 984
rect 6166 202 6172 984
rect 6108 198 6172 202
rect 6266 980 6330 986
rect 6266 202 6272 980
rect 6324 202 6330 980
rect 5957 192 6003 196
rect 6115 192 6161 198
rect 6266 196 6330 202
rect 6424 984 6488 988
rect 6589 986 6635 992
rect 6747 988 6793 992
rect 6424 202 6430 984
rect 6482 202 6488 984
rect 6424 198 6488 202
rect 6582 980 6646 986
rect 6582 202 6588 980
rect 6640 202 6646 980
rect 6273 192 6319 196
rect 6431 192 6477 198
rect 6582 196 6646 202
rect 6740 984 6804 988
rect 6905 986 6951 992
rect 7063 988 7109 992
rect 6740 202 6746 984
rect 6798 202 6804 984
rect 6740 198 6804 202
rect 6898 980 6962 986
rect 6898 202 6904 980
rect 6956 202 6962 980
rect 6589 192 6635 196
rect 6747 192 6793 198
rect 6898 196 6962 202
rect 7056 984 7120 988
rect 7221 986 7267 992
rect 7379 988 7425 992
rect 7056 202 7062 984
rect 7114 202 7120 984
rect 7056 198 7120 202
rect 7214 980 7278 986
rect 7214 202 7220 980
rect 7272 202 7278 980
rect 6905 192 6951 196
rect 7063 192 7109 198
rect 7214 196 7278 202
rect 7372 984 7436 988
rect 7537 986 7583 992
rect 7695 988 7741 992
rect 7372 202 7378 984
rect 7430 202 7436 984
rect 7372 198 7436 202
rect 7530 980 7594 986
rect 7530 202 7536 980
rect 7588 202 7594 980
rect 7221 192 7267 196
rect 7379 192 7425 198
rect 7530 196 7594 202
rect 7688 984 7752 988
rect 7853 986 7899 992
rect 8011 988 8057 992
rect 7688 202 7694 984
rect 7746 202 7752 984
rect 7688 198 7752 202
rect 7846 980 7910 986
rect 7846 202 7852 980
rect 7904 202 7910 980
rect 7537 192 7583 196
rect 7695 192 7741 198
rect 7846 196 7910 202
rect 8004 984 8068 988
rect 8169 986 8215 992
rect 8327 988 8373 992
rect 8004 202 8010 984
rect 8062 202 8068 984
rect 8004 198 8068 202
rect 8162 980 8226 986
rect 8162 202 8168 980
rect 8220 202 8226 980
rect 7853 192 7899 196
rect 8011 192 8057 198
rect 8162 196 8226 202
rect 8320 984 8384 988
rect 8485 986 8531 992
rect 8643 988 8689 992
rect 8320 202 8326 984
rect 8378 202 8384 984
rect 8320 198 8384 202
rect 8478 980 8542 986
rect 8478 202 8484 980
rect 8536 202 8542 980
rect 8169 192 8215 196
rect 8327 192 8373 198
rect 8478 196 8542 202
rect 8636 984 8700 988
rect 8801 986 8847 992
rect 8959 988 9005 992
rect 8636 202 8642 984
rect 8694 202 8700 984
rect 8636 198 8700 202
rect 8794 980 8858 986
rect 8794 202 8800 980
rect 8852 202 8858 980
rect 8485 192 8531 196
rect 8643 192 8689 198
rect 8794 196 8858 202
rect 8952 984 9016 988
rect 9117 986 9163 992
rect 9275 988 9321 992
rect 8952 202 8958 984
rect 9010 202 9016 984
rect 8952 198 9016 202
rect 9110 980 9174 986
rect 9110 202 9116 980
rect 9168 202 9174 980
rect 8801 192 8847 196
rect 8959 192 9005 198
rect 9110 196 9174 202
rect 9268 984 9332 988
rect 9433 986 9479 992
rect 9591 988 9637 992
rect 9268 202 9274 984
rect 9326 202 9332 984
rect 9268 198 9332 202
rect 9426 980 9490 986
rect 9426 202 9432 980
rect 9484 202 9490 980
rect 9117 192 9163 196
rect 9275 192 9321 198
rect 9426 196 9490 202
rect 9584 984 9648 988
rect 9749 986 9795 992
rect 9907 988 9953 992
rect 9584 202 9590 984
rect 9642 202 9648 984
rect 9584 198 9648 202
rect 9742 980 9806 986
rect 9742 202 9748 980
rect 9800 202 9806 980
rect 9433 192 9479 196
rect 9591 192 9637 198
rect 9742 196 9806 202
rect 9900 984 9964 988
rect 10065 986 10111 992
rect 10223 988 10269 992
rect 9900 202 9906 984
rect 9958 202 9964 984
rect 9900 198 9964 202
rect 10058 980 10122 986
rect 10058 202 10064 980
rect 10116 202 10122 980
rect 9749 192 9795 196
rect 9907 192 9953 198
rect 10058 196 10122 202
rect 10216 984 10280 988
rect 10381 986 10427 992
rect 10539 988 10585 992
rect 10216 202 10222 984
rect 10274 202 10280 984
rect 10216 198 10280 202
rect 10374 980 10438 986
rect 10374 202 10380 980
rect 10432 202 10438 980
rect 10065 192 10111 196
rect 10223 192 10269 198
rect 10374 196 10438 202
rect 10532 984 10596 988
rect 10697 986 10743 992
rect 10855 988 10901 992
rect 10532 202 10538 984
rect 10590 202 10596 984
rect 10532 198 10596 202
rect 10690 980 10754 986
rect 10690 202 10696 980
rect 10748 202 10754 980
rect 10381 192 10427 196
rect 10539 192 10585 198
rect 10690 196 10754 202
rect 10848 984 10912 988
rect 11013 986 11059 992
rect 11171 988 11217 992
rect 10848 202 10854 984
rect 10906 202 10912 984
rect 10848 198 10912 202
rect 11006 980 11070 986
rect 11006 202 11012 980
rect 11064 202 11070 980
rect 10697 192 10743 196
rect 10855 192 10901 198
rect 11006 196 11070 202
rect 11164 984 11228 988
rect 11329 986 11375 992
rect 11487 988 11533 992
rect 11164 202 11170 984
rect 11222 202 11228 984
rect 11164 198 11228 202
rect 11322 980 11386 986
rect 11322 202 11328 980
rect 11380 202 11386 980
rect 11013 192 11059 196
rect 11171 192 11217 198
rect 11322 196 11386 202
rect 11480 984 11544 988
rect 11645 986 11691 992
rect 11803 988 11849 992
rect 11480 202 11486 984
rect 11538 202 11544 984
rect 11480 198 11544 202
rect 11638 980 11702 986
rect 11638 202 11644 980
rect 11696 202 11702 980
rect 11329 192 11375 196
rect 11487 192 11533 198
rect 11638 196 11702 202
rect 11796 984 11860 988
rect 11961 986 12007 992
rect 12119 988 12165 992
rect 11796 202 11802 984
rect 11854 202 11860 984
rect 11796 198 11860 202
rect 11954 980 12018 986
rect 11954 202 11960 980
rect 12012 202 12018 980
rect 11645 192 11691 196
rect 11803 192 11849 198
rect 11954 196 12018 202
rect 12112 984 12176 988
rect 12277 986 12323 992
rect 12435 988 12481 992
rect 12112 202 12118 984
rect 12170 202 12176 984
rect 12112 198 12176 202
rect 12270 980 12334 986
rect 12270 202 12276 980
rect 12328 202 12334 980
rect 11961 192 12007 196
rect 12119 192 12165 198
rect 12270 196 12334 202
rect 12428 984 12492 988
rect 12593 986 12639 992
rect 12745 988 12791 992
rect 12428 202 12434 984
rect 12486 202 12492 984
rect 12428 198 12492 202
rect 12586 980 12650 986
rect 12586 202 12592 980
rect 12644 202 12650 980
rect 12277 192 12323 196
rect 12435 192 12481 198
rect 12586 196 12650 202
rect 12738 984 12802 988
rect 12738 202 12744 984
rect 12796 202 12802 984
rect 12738 198 12802 202
rect 12593 192 12639 196
rect 12745 192 12791 198
rect 12830 160 12864 1024
rect 42 114 12864 160
rect 12892 1932 12950 1972
rect 254 26 330 32
rect 254 16 260 26
rect 324 16 330 26
rect 570 26 646 32
rect 570 16 576 26
rect 640 16 646 26
rect 886 26 962 32
rect 886 16 892 26
rect 956 16 962 26
rect 1202 26 1278 32
rect 1202 16 1208 26
rect 1272 16 1278 26
rect 1518 26 1594 32
rect 1518 16 1524 26
rect 1588 16 1594 26
rect 1834 26 1910 32
rect 1834 16 1840 26
rect 1904 16 1910 26
rect 2150 26 2226 32
rect 2150 16 2156 26
rect 2220 16 2226 26
rect 2466 26 2542 32
rect 2466 16 2472 26
rect 2536 16 2542 26
rect 2782 26 2858 32
rect 2782 16 2788 26
rect 2852 16 2858 26
rect 3098 26 3174 32
rect 3098 16 3104 26
rect 3168 16 3174 26
rect 3414 26 3490 32
rect 3414 16 3420 26
rect 3484 16 3490 26
rect 3730 26 3806 32
rect 3730 16 3736 26
rect 3800 16 3806 26
rect 4046 26 4122 32
rect 4046 16 4052 26
rect 4116 16 4122 26
rect 4362 26 4438 32
rect 4362 16 4368 26
rect 4432 16 4438 26
rect 4678 26 4754 32
rect 4678 16 4684 26
rect 4748 16 4754 26
rect 4994 26 5070 32
rect 4994 16 5000 26
rect 5064 16 5070 26
rect 5310 26 5386 32
rect 5310 16 5316 26
rect 5380 16 5386 26
rect 5626 26 5702 32
rect 5626 16 5632 26
rect 5696 16 5702 26
rect 5942 26 6018 32
rect 5942 16 5948 26
rect 6012 16 6018 26
rect 6258 26 6334 32
rect 6258 16 6264 26
rect 6328 16 6334 26
rect 6574 26 6650 32
rect 6574 16 6580 26
rect 6644 16 6650 26
rect 6890 26 6966 32
rect 6890 16 6896 26
rect 6960 16 6966 26
rect 7206 26 7282 32
rect 7206 16 7212 26
rect 7276 16 7282 26
rect 7522 26 7598 32
rect 7522 16 7528 26
rect 7592 16 7598 26
rect 7838 26 7914 32
rect 7838 16 7844 26
rect 7908 16 7914 26
rect 8154 26 8230 32
rect 8154 16 8160 26
rect 8224 16 8230 26
rect 8470 26 8546 32
rect 8470 16 8476 26
rect 8540 16 8546 26
rect 8786 26 8862 32
rect 8786 16 8792 26
rect 8856 16 8862 26
rect 9102 26 9178 32
rect 9102 16 9108 26
rect 9172 16 9178 26
rect 9418 26 9494 32
rect 9418 16 9424 26
rect 9488 16 9494 26
rect 9734 26 9810 32
rect 9734 16 9740 26
rect 9804 16 9810 26
rect 10050 26 10126 32
rect 10050 16 10056 26
rect 10120 16 10126 26
rect 10366 26 10442 32
rect 10366 16 10372 26
rect 10436 16 10442 26
rect 10682 26 10758 32
rect 10682 16 10688 26
rect 10752 16 10758 26
rect 10998 26 11074 32
rect 10998 16 11004 26
rect 11068 16 11074 26
rect 11314 26 11390 32
rect 11314 16 11320 26
rect 11384 16 11390 26
rect 11630 26 11706 32
rect 11630 16 11636 26
rect 11700 16 11706 26
rect 11946 26 12022 32
rect 11946 16 11952 26
rect 12016 16 12022 26
rect 12262 26 12338 32
rect 12262 16 12268 26
rect 12332 16 12338 26
rect 12578 26 12654 32
rect 12578 16 12584 26
rect 12648 16 12654 26
rect 12892 16 12904 1932
rect 2 -6 260 16
rect -44 -18 260 -6
rect 324 -18 576 16
rect 640 -18 892 16
rect 956 -18 1208 16
rect 1272 -18 1524 16
rect 1588 -18 1840 16
rect 1904 -18 2156 16
rect 2220 -18 2472 16
rect 2536 -18 2788 16
rect 2852 -18 3104 16
rect 3168 -18 3420 16
rect 3484 -18 3736 16
rect 3800 -18 4052 16
rect 4116 -18 4368 16
rect 4432 -18 4684 16
rect 4748 -18 5000 16
rect 5064 -18 5316 16
rect 5380 -18 5632 16
rect 5696 -18 5948 16
rect 6012 -18 6264 16
rect 6328 -18 6580 16
rect 6644 -18 6896 16
rect 6960 -18 7212 16
rect 7276 -18 7528 16
rect 7592 -18 7844 16
rect 7908 -18 8160 16
rect 8224 -18 8476 16
rect 8540 -18 8792 16
rect 8856 -18 9108 16
rect 9172 -18 9424 16
rect 9488 -18 9740 16
rect 9804 -18 10056 16
rect 10120 -18 10372 16
rect 10436 -18 10688 16
rect 10752 -18 11004 16
rect 11068 -18 11320 16
rect 11384 -18 11636 16
rect 11700 -18 11952 16
rect 12016 -18 12268 16
rect 12332 -18 12584 16
rect 12648 -6 12904 16
rect 12938 -6 12950 1932
rect 12648 -18 12950 -6
rect 254 -28 260 -18
rect 324 -28 330 -18
rect 254 -34 330 -28
rect 570 -28 576 -18
rect 640 -28 646 -18
rect 570 -34 646 -28
rect 886 -28 892 -18
rect 956 -28 962 -18
rect 886 -34 962 -28
rect 1202 -28 1208 -18
rect 1272 -28 1278 -18
rect 1202 -34 1278 -28
rect 1518 -28 1524 -18
rect 1588 -28 1594 -18
rect 1518 -34 1594 -28
rect 1834 -28 1840 -18
rect 1904 -28 1910 -18
rect 1834 -34 1910 -28
rect 2150 -28 2156 -18
rect 2220 -28 2226 -18
rect 2150 -34 2226 -28
rect 2466 -28 2472 -18
rect 2536 -28 2542 -18
rect 2466 -34 2542 -28
rect 2782 -28 2788 -18
rect 2852 -28 2858 -18
rect 2782 -34 2858 -28
rect 3098 -28 3104 -18
rect 3168 -28 3174 -18
rect 3098 -34 3174 -28
rect 3414 -28 3420 -18
rect 3484 -28 3490 -18
rect 3414 -34 3490 -28
rect 3730 -28 3736 -18
rect 3800 -28 3806 -18
rect 3730 -34 3806 -28
rect 4046 -28 4052 -18
rect 4116 -28 4122 -18
rect 4046 -34 4122 -28
rect 4362 -28 4368 -18
rect 4432 -28 4438 -18
rect 4362 -34 4438 -28
rect 4678 -28 4684 -18
rect 4748 -28 4754 -18
rect 4678 -34 4754 -28
rect 4994 -28 5000 -18
rect 5064 -28 5070 -18
rect 4994 -34 5070 -28
rect 5310 -28 5316 -18
rect 5380 -28 5386 -18
rect 5310 -34 5386 -28
rect 5626 -28 5632 -18
rect 5696 -28 5702 -18
rect 5626 -34 5702 -28
rect 5942 -28 5948 -18
rect 6012 -28 6018 -18
rect 5942 -34 6018 -28
rect 6258 -28 6264 -18
rect 6328 -28 6334 -18
rect 6258 -34 6334 -28
rect 6574 -28 6580 -18
rect 6644 -28 6650 -18
rect 6574 -34 6650 -28
rect 6890 -28 6896 -18
rect 6960 -28 6966 -18
rect 6890 -34 6966 -28
rect 7206 -28 7212 -18
rect 7276 -28 7282 -18
rect 7206 -34 7282 -28
rect 7522 -28 7528 -18
rect 7592 -28 7598 -18
rect 7522 -34 7598 -28
rect 7838 -28 7844 -18
rect 7908 -28 7914 -18
rect 7838 -34 7914 -28
rect 8154 -28 8160 -18
rect 8224 -28 8230 -18
rect 8154 -34 8230 -28
rect 8470 -28 8476 -18
rect 8540 -28 8546 -18
rect 8470 -34 8546 -28
rect 8786 -28 8792 -18
rect 8856 -28 8862 -18
rect 8786 -34 8862 -28
rect 9102 -28 9108 -18
rect 9172 -28 9178 -18
rect 9102 -34 9178 -28
rect 9418 -28 9424 -18
rect 9488 -28 9494 -18
rect 9418 -34 9494 -28
rect 9734 -28 9740 -18
rect 9804 -28 9810 -18
rect 9734 -34 9810 -28
rect 10050 -28 10056 -18
rect 10120 -28 10126 -18
rect 10050 -34 10126 -28
rect 10366 -28 10372 -18
rect 10436 -28 10442 -18
rect 10366 -34 10442 -28
rect 10682 -28 10688 -18
rect 10752 -28 10758 -18
rect 10682 -34 10758 -28
rect 10998 -28 11004 -18
rect 11068 -28 11074 -18
rect 10998 -34 11074 -28
rect 11314 -28 11320 -18
rect 11384 -28 11390 -18
rect 11314 -34 11390 -28
rect 11630 -28 11636 -18
rect 11700 -28 11706 -18
rect 11630 -34 11706 -28
rect 11946 -28 11952 -18
rect 12016 -28 12022 -18
rect 11946 -34 12022 -28
rect 12262 -28 12268 -18
rect 12332 -28 12338 -18
rect 12262 -34 12338 -28
rect 12578 -28 12584 -18
rect 12648 -28 12654 -18
rect 12578 -34 12654 -28
<< via1 >>
rect 260 4842 324 4852
rect 576 4842 640 4852
rect 892 4842 956 4852
rect 1208 4842 1272 4852
rect 1524 4842 1588 4852
rect 1840 4842 1904 4852
rect 2156 4842 2220 4852
rect 2472 4842 2536 4852
rect 2788 4842 2852 4852
rect 3104 4842 3168 4852
rect 3420 4842 3484 4852
rect 3736 4842 3800 4852
rect 4052 4842 4116 4852
rect 4368 4842 4432 4852
rect 4684 4842 4748 4852
rect 5000 4842 5064 4852
rect 5316 4842 5380 4852
rect 5632 4842 5696 4852
rect 5948 4842 6012 4852
rect 6264 4842 6328 4852
rect 6580 4842 6644 4852
rect 6896 4842 6960 4852
rect 7212 4842 7276 4852
rect 7528 4842 7592 4852
rect 7844 4842 7908 4852
rect 8160 4842 8224 4852
rect 8476 4842 8540 4852
rect 8792 4842 8856 4852
rect 9108 4842 9172 4852
rect 9424 4842 9488 4852
rect 9740 4842 9804 4852
rect 10056 4842 10120 4852
rect 10372 4842 10436 4852
rect 10688 4842 10752 4852
rect 11004 4842 11068 4852
rect 11320 4842 11384 4852
rect 11636 4842 11700 4852
rect 11952 4842 12016 4852
rect 12268 4842 12332 4852
rect 12584 4842 12648 4852
rect 260 4808 274 4842
rect 274 4808 310 4842
rect 310 4808 324 4842
rect 576 4808 590 4842
rect 590 4808 626 4842
rect 626 4808 640 4842
rect 892 4808 906 4842
rect 906 4808 942 4842
rect 942 4808 956 4842
rect 1208 4808 1222 4842
rect 1222 4808 1258 4842
rect 1258 4808 1272 4842
rect 1524 4808 1538 4842
rect 1538 4808 1574 4842
rect 1574 4808 1588 4842
rect 1840 4808 1854 4842
rect 1854 4808 1890 4842
rect 1890 4808 1904 4842
rect 2156 4808 2170 4842
rect 2170 4808 2206 4842
rect 2206 4808 2220 4842
rect 2472 4808 2486 4842
rect 2486 4808 2522 4842
rect 2522 4808 2536 4842
rect 2788 4808 2802 4842
rect 2802 4808 2838 4842
rect 2838 4808 2852 4842
rect 3104 4808 3118 4842
rect 3118 4808 3154 4842
rect 3154 4808 3168 4842
rect 3420 4808 3434 4842
rect 3434 4808 3470 4842
rect 3470 4808 3484 4842
rect 3736 4808 3750 4842
rect 3750 4808 3786 4842
rect 3786 4808 3800 4842
rect 4052 4808 4066 4842
rect 4066 4808 4102 4842
rect 4102 4808 4116 4842
rect 4368 4808 4382 4842
rect 4382 4808 4418 4842
rect 4418 4808 4432 4842
rect 4684 4808 4698 4842
rect 4698 4808 4734 4842
rect 4734 4808 4748 4842
rect 5000 4808 5014 4842
rect 5014 4808 5050 4842
rect 5050 4808 5064 4842
rect 5316 4808 5330 4842
rect 5330 4808 5366 4842
rect 5366 4808 5380 4842
rect 5632 4808 5646 4842
rect 5646 4808 5682 4842
rect 5682 4808 5696 4842
rect 5948 4808 5962 4842
rect 5962 4808 5998 4842
rect 5998 4808 6012 4842
rect 6264 4808 6278 4842
rect 6278 4808 6314 4842
rect 6314 4808 6328 4842
rect 6580 4808 6594 4842
rect 6594 4808 6630 4842
rect 6630 4808 6644 4842
rect 6896 4808 6910 4842
rect 6910 4808 6946 4842
rect 6946 4808 6960 4842
rect 7212 4808 7226 4842
rect 7226 4808 7262 4842
rect 7262 4808 7276 4842
rect 7528 4808 7542 4842
rect 7542 4808 7578 4842
rect 7578 4808 7592 4842
rect 7844 4808 7858 4842
rect 7858 4808 7894 4842
rect 7894 4808 7908 4842
rect 8160 4808 8174 4842
rect 8174 4808 8210 4842
rect 8210 4808 8224 4842
rect 8476 4808 8490 4842
rect 8490 4808 8526 4842
rect 8526 4808 8540 4842
rect 8792 4808 8806 4842
rect 8806 4808 8842 4842
rect 8842 4808 8856 4842
rect 9108 4808 9122 4842
rect 9122 4808 9158 4842
rect 9158 4808 9172 4842
rect 9424 4808 9438 4842
rect 9438 4808 9474 4842
rect 9474 4808 9488 4842
rect 9740 4808 9754 4842
rect 9754 4808 9790 4842
rect 9790 4808 9804 4842
rect 10056 4808 10070 4842
rect 10070 4808 10106 4842
rect 10106 4808 10120 4842
rect 10372 4808 10386 4842
rect 10386 4808 10422 4842
rect 10422 4808 10436 4842
rect 10688 4808 10702 4842
rect 10702 4808 10738 4842
rect 10738 4808 10752 4842
rect 11004 4808 11018 4842
rect 11018 4808 11054 4842
rect 11054 4808 11068 4842
rect 11320 4808 11334 4842
rect 11334 4808 11370 4842
rect 11370 4808 11384 4842
rect 11636 4808 11650 4842
rect 11650 4808 11686 4842
rect 11686 4808 11700 4842
rect 11952 4808 11966 4842
rect 11966 4808 12002 4842
rect 12002 4808 12016 4842
rect 12268 4808 12282 4842
rect 12282 4808 12318 4842
rect 12318 4808 12332 4842
rect 12584 4808 12598 4842
rect 12598 4808 12634 4842
rect 12634 4808 12648 4842
rect 260 4798 324 4808
rect 576 4798 640 4808
rect 892 4798 956 4808
rect 1208 4798 1272 4808
rect 1524 4798 1588 4808
rect 1840 4798 1904 4808
rect 2156 4798 2220 4808
rect 2472 4798 2536 4808
rect 2788 4798 2852 4808
rect 3104 4798 3168 4808
rect 3420 4798 3484 4808
rect 3736 4798 3800 4808
rect 4052 4798 4116 4808
rect 4368 4798 4432 4808
rect 4684 4798 4748 4808
rect 5000 4798 5064 4808
rect 5316 4798 5380 4808
rect 5632 4798 5696 4808
rect 5948 4798 6012 4808
rect 6264 4798 6328 4808
rect 6580 4798 6644 4808
rect 6896 4798 6960 4808
rect 7212 4798 7276 4808
rect 7528 4798 7592 4808
rect 7844 4798 7908 4808
rect 8160 4798 8224 4808
rect 8476 4798 8540 4808
rect 8792 4798 8856 4808
rect 9108 4798 9172 4808
rect 9424 4798 9488 4808
rect 9740 4798 9804 4808
rect 10056 4798 10120 4808
rect 10372 4798 10436 4808
rect 10688 4798 10752 4808
rect 11004 4798 11068 4808
rect 11320 4798 11384 4808
rect 11636 4798 11700 4808
rect 11952 4798 12016 4808
rect 12268 4798 12332 4808
rect 12584 4798 12648 4808
rect 110 3844 162 4622
rect 268 3840 320 4622
rect 426 3844 478 4622
rect 584 3840 636 4622
rect 742 3844 794 4622
rect 900 3840 952 4622
rect 1058 3844 1110 4622
rect 1216 3840 1268 4622
rect 1374 3844 1426 4622
rect 1532 3840 1584 4622
rect 1690 3844 1742 4622
rect 1848 3840 1900 4622
rect 2006 3844 2058 4622
rect 2164 3840 2216 4622
rect 2322 3844 2374 4622
rect 2480 3840 2532 4622
rect 2638 3844 2690 4622
rect 2796 3840 2848 4622
rect 2954 3844 3006 4622
rect 3112 3840 3164 4622
rect 3270 3844 3322 4622
rect 3428 3840 3480 4622
rect 3586 3844 3638 4622
rect 3744 3840 3796 4622
rect 3902 3844 3954 4622
rect 4060 3840 4112 4622
rect 4218 3844 4270 4622
rect 4376 3840 4428 4622
rect 4534 3844 4586 4622
rect 4692 3840 4744 4622
rect 4850 3844 4902 4622
rect 5008 3840 5060 4622
rect 5166 3844 5218 4622
rect 5324 3840 5376 4622
rect 5482 3844 5534 4622
rect 5640 3840 5692 4622
rect 5798 3844 5850 4622
rect 5956 3840 6008 4622
rect 6114 3844 6166 4622
rect 6272 3840 6324 4622
rect 6430 3844 6482 4622
rect 6588 3840 6640 4622
rect 6746 3844 6798 4622
rect 6904 3840 6956 4622
rect 7062 3844 7114 4622
rect 7220 3840 7272 4622
rect 7378 3844 7430 4622
rect 7536 3840 7588 4622
rect 7694 3844 7746 4622
rect 7852 3840 7904 4622
rect 8010 3844 8062 4622
rect 8168 3840 8220 4622
rect 8326 3844 8378 4622
rect 8484 3840 8536 4622
rect 8642 3844 8694 4622
rect 8800 3840 8852 4622
rect 8958 3844 9010 4622
rect 9116 3840 9168 4622
rect 9274 3844 9326 4622
rect 9432 3840 9484 4622
rect 9590 3844 9642 4622
rect 9748 3840 9800 4622
rect 9906 3844 9958 4622
rect 10064 3840 10116 4622
rect 10222 3844 10274 4622
rect 10380 3840 10432 4622
rect 10538 3844 10590 4622
rect 10696 3840 10748 4622
rect 10854 3844 10906 4622
rect 11012 3840 11064 4622
rect 11170 3844 11222 4622
rect 11328 3840 11380 4622
rect 11486 3844 11538 4622
rect 11644 3840 11696 4622
rect 11802 3844 11854 4622
rect 11960 3840 12012 4622
rect 12118 3844 12170 4622
rect 12276 3840 12328 4622
rect 12434 3844 12486 4622
rect 12592 3840 12644 4622
rect 12744 3844 12796 4622
rect 110 2932 162 3714
rect 268 2930 320 3712
rect 426 2932 478 3714
rect 584 2930 636 3712
rect 742 2932 794 3714
rect 900 2930 952 3712
rect 1058 2932 1110 3714
rect 1216 2930 1268 3712
rect 1374 2932 1426 3714
rect 1532 2930 1584 3712
rect 1690 2932 1742 3714
rect 1848 2930 1900 3712
rect 2006 2932 2058 3714
rect 2164 2930 2216 3712
rect 2322 2932 2374 3714
rect 2480 2930 2532 3712
rect 2638 2932 2690 3714
rect 2796 2930 2848 3712
rect 2954 2932 3006 3714
rect 3112 2930 3164 3712
rect 3270 2932 3322 3714
rect 3428 2930 3480 3712
rect 3586 2932 3638 3714
rect 3744 2930 3796 3712
rect 3902 2932 3954 3714
rect 4060 2930 4112 3712
rect 4218 2932 4270 3714
rect 4376 2930 4428 3712
rect 4534 2932 4586 3714
rect 4692 2930 4744 3712
rect 4850 2932 4902 3714
rect 5008 2930 5060 3712
rect 5166 2932 5218 3714
rect 5324 2930 5376 3712
rect 5482 2932 5534 3714
rect 5640 2930 5692 3712
rect 5798 2932 5850 3714
rect 5956 2930 6008 3712
rect 6114 2932 6166 3714
rect 6272 2930 6324 3712
rect 6430 2932 6482 3714
rect 6588 2930 6640 3712
rect 6746 2932 6798 3714
rect 6904 2930 6956 3712
rect 7062 2932 7114 3714
rect 7220 2930 7272 3712
rect 7378 2932 7430 3714
rect 7536 2930 7588 3712
rect 7694 2932 7746 3714
rect 7852 2930 7904 3712
rect 8010 2932 8062 3714
rect 8168 2930 8220 3712
rect 8326 2932 8378 3714
rect 8484 2930 8536 3712
rect 8642 2932 8694 3714
rect 8800 2930 8852 3712
rect 8958 2932 9010 3714
rect 9116 2930 9168 3712
rect 9274 2932 9326 3714
rect 9432 2930 9484 3712
rect 9590 2932 9642 3714
rect 9748 2930 9800 3712
rect 9906 2932 9958 3714
rect 10064 2930 10116 3712
rect 10222 2932 10274 3714
rect 10380 2930 10432 3712
rect 10538 2932 10590 3714
rect 10696 2930 10748 3712
rect 10854 2932 10906 3714
rect 11012 2930 11064 3712
rect 11170 2932 11222 3714
rect 11328 2930 11380 3712
rect 11486 2932 11538 3714
rect 11644 2930 11696 3712
rect 11802 2932 11854 3714
rect 11960 2930 12012 3712
rect 12118 2932 12170 3714
rect 12276 2930 12328 3712
rect 12434 2932 12486 3714
rect 12592 2930 12644 3712
rect 12744 2932 12796 3714
rect 110 2022 162 2804
rect 268 2020 320 2802
rect 426 2022 478 2804
rect 584 2020 636 2802
rect 742 2022 794 2804
rect 900 2020 952 2802
rect 1058 2022 1110 2804
rect 1216 2020 1268 2802
rect 1374 2022 1426 2804
rect 1532 2020 1584 2802
rect 1690 2022 1742 2804
rect 1848 2020 1900 2802
rect 2006 2022 2058 2804
rect 2164 2020 2216 2802
rect 2322 2022 2374 2804
rect 2480 2020 2532 2802
rect 2638 2022 2690 2804
rect 2796 2020 2848 2802
rect 2954 2022 3006 2804
rect 3112 2020 3164 2802
rect 3270 2022 3322 2804
rect 3428 2020 3480 2802
rect 3586 2022 3638 2804
rect 3744 2020 3796 2802
rect 3902 2022 3954 2804
rect 4060 2020 4112 2802
rect 4218 2022 4270 2804
rect 4376 2020 4428 2802
rect 4534 2022 4586 2804
rect 4692 2020 4744 2802
rect 4850 2022 4902 2804
rect 5008 2020 5060 2802
rect 5166 2022 5218 2804
rect 5324 2020 5376 2802
rect 5482 2022 5534 2804
rect 5640 2020 5692 2802
rect 5798 2022 5850 2804
rect 5956 2020 6008 2802
rect 6114 2022 6166 2804
rect 6272 2020 6324 2802
rect 6430 2022 6482 2804
rect 6588 2020 6640 2802
rect 6746 2022 6798 2804
rect 6904 2020 6956 2802
rect 7062 2022 7114 2804
rect 7220 2020 7272 2802
rect 7378 2022 7430 2804
rect 7536 2020 7588 2802
rect 7694 2022 7746 2804
rect 7852 2020 7904 2802
rect 8010 2022 8062 2804
rect 8168 2020 8220 2802
rect 8326 2022 8378 2804
rect 8484 2020 8536 2802
rect 8642 2022 8694 2804
rect 8800 2020 8852 2802
rect 8958 2022 9010 2804
rect 9116 2020 9168 2802
rect 9274 2022 9326 2804
rect 9432 2020 9484 2802
rect 9590 2022 9642 2804
rect 9748 2020 9800 2802
rect 9906 2022 9958 2804
rect 10064 2020 10116 2802
rect 10222 2022 10274 2804
rect 10380 2020 10432 2802
rect 10538 2022 10590 2804
rect 10696 2020 10748 2802
rect 10854 2022 10906 2804
rect 11012 2020 11064 2802
rect 11170 2022 11222 2804
rect 11328 2020 11380 2802
rect 11486 2022 11538 2804
rect 11644 2020 11696 2802
rect 11802 2022 11854 2804
rect 11960 2020 12012 2802
rect 12118 2022 12170 2804
rect 12276 2020 12328 2802
rect 12434 2022 12486 2804
rect 12592 2020 12644 2802
rect 12744 2022 12796 2804
rect 110 1112 162 1894
rect 268 1110 320 1892
rect 426 1112 478 1894
rect 584 1110 636 1892
rect 742 1112 794 1894
rect 900 1110 952 1892
rect 1058 1112 1110 1894
rect 1216 1110 1268 1892
rect 1374 1112 1426 1894
rect 1532 1110 1584 1892
rect 1690 1112 1742 1894
rect 1848 1110 1900 1892
rect 2006 1112 2058 1894
rect 2164 1110 2216 1892
rect 2322 1112 2374 1894
rect 2480 1110 2532 1892
rect 2638 1112 2690 1894
rect 2796 1110 2848 1892
rect 2954 1112 3006 1894
rect 3112 1110 3164 1892
rect 3270 1112 3322 1894
rect 3428 1110 3480 1892
rect 3586 1112 3638 1894
rect 3744 1110 3796 1892
rect 3902 1112 3954 1894
rect 4060 1110 4112 1892
rect 4218 1112 4270 1894
rect 4376 1110 4428 1892
rect 4534 1112 4586 1894
rect 4692 1110 4744 1892
rect 4850 1112 4902 1894
rect 5008 1110 5060 1892
rect 5166 1112 5218 1894
rect 5324 1110 5376 1892
rect 5482 1112 5534 1894
rect 5640 1110 5692 1892
rect 5798 1112 5850 1894
rect 5956 1110 6008 1892
rect 6114 1112 6166 1894
rect 6272 1110 6324 1892
rect 6430 1112 6482 1894
rect 6588 1110 6640 1892
rect 6746 1112 6798 1894
rect 6904 1110 6956 1892
rect 7062 1112 7114 1894
rect 7220 1110 7272 1892
rect 7378 1112 7430 1894
rect 7536 1110 7588 1892
rect 7694 1112 7746 1894
rect 7852 1110 7904 1892
rect 8010 1112 8062 1894
rect 8168 1110 8220 1892
rect 8326 1112 8378 1894
rect 8484 1110 8536 1892
rect 8642 1112 8694 1894
rect 8800 1110 8852 1892
rect 8958 1112 9010 1894
rect 9116 1110 9168 1892
rect 9274 1112 9326 1894
rect 9432 1110 9484 1892
rect 9590 1112 9642 1894
rect 9748 1110 9800 1892
rect 9906 1112 9958 1894
rect 10064 1110 10116 1892
rect 10222 1112 10274 1894
rect 10380 1110 10432 1892
rect 10538 1112 10590 1894
rect 10696 1110 10748 1892
rect 10854 1112 10906 1894
rect 11012 1110 11064 1892
rect 11170 1112 11222 1894
rect 11328 1110 11380 1892
rect 11486 1112 11538 1894
rect 11644 1110 11696 1892
rect 11802 1112 11854 1894
rect 11960 1110 12012 1892
rect 12118 1112 12170 1894
rect 12276 1110 12328 1892
rect 12434 1112 12486 1894
rect 12592 1110 12644 1892
rect 12744 1112 12796 1894
rect 110 202 162 984
rect 268 202 320 980
rect 426 202 478 984
rect 584 202 636 980
rect 742 202 794 984
rect 900 202 952 980
rect 1058 202 1110 984
rect 1216 202 1268 980
rect 1374 202 1426 984
rect 1532 202 1584 980
rect 1690 202 1742 984
rect 1848 202 1900 980
rect 2006 202 2058 984
rect 2164 202 2216 980
rect 2322 202 2374 984
rect 2480 202 2532 980
rect 2638 202 2690 984
rect 2796 202 2848 980
rect 2954 202 3006 984
rect 3112 202 3164 980
rect 3270 202 3322 984
rect 3428 202 3480 980
rect 3586 202 3638 984
rect 3744 202 3796 980
rect 3902 202 3954 984
rect 4060 202 4112 980
rect 4218 202 4270 984
rect 4376 202 4428 980
rect 4534 202 4586 984
rect 4692 202 4744 980
rect 4850 202 4902 984
rect 5008 202 5060 980
rect 5166 202 5218 984
rect 5324 202 5376 980
rect 5482 202 5534 984
rect 5640 202 5692 980
rect 5798 202 5850 984
rect 5956 202 6008 980
rect 6114 202 6166 984
rect 6272 202 6324 980
rect 6430 202 6482 984
rect 6588 202 6640 980
rect 6746 202 6798 984
rect 6904 202 6956 980
rect 7062 202 7114 984
rect 7220 202 7272 980
rect 7378 202 7430 984
rect 7536 202 7588 980
rect 7694 202 7746 984
rect 7852 202 7904 980
rect 8010 202 8062 984
rect 8168 202 8220 980
rect 8326 202 8378 984
rect 8484 202 8536 980
rect 8642 202 8694 984
rect 8800 202 8852 980
rect 8958 202 9010 984
rect 9116 202 9168 980
rect 9274 202 9326 984
rect 9432 202 9484 980
rect 9590 202 9642 984
rect 9748 202 9800 980
rect 9906 202 9958 984
rect 10064 202 10116 980
rect 10222 202 10274 984
rect 10380 202 10432 980
rect 10538 202 10590 984
rect 10696 202 10748 980
rect 10854 202 10906 984
rect 11012 202 11064 980
rect 11170 202 11222 984
rect 11328 202 11380 980
rect 11486 202 11538 984
rect 11644 202 11696 980
rect 11802 202 11854 984
rect 11960 202 12012 980
rect 12118 202 12170 984
rect 12276 202 12328 980
rect 12434 202 12486 984
rect 12592 202 12644 980
rect 12744 202 12796 984
rect 260 16 324 26
rect 576 16 640 26
rect 892 16 956 26
rect 1208 16 1272 26
rect 1524 16 1588 26
rect 1840 16 1904 26
rect 2156 16 2220 26
rect 2472 16 2536 26
rect 2788 16 2852 26
rect 3104 16 3168 26
rect 3420 16 3484 26
rect 3736 16 3800 26
rect 4052 16 4116 26
rect 4368 16 4432 26
rect 4684 16 4748 26
rect 5000 16 5064 26
rect 5316 16 5380 26
rect 5632 16 5696 26
rect 5948 16 6012 26
rect 6264 16 6328 26
rect 6580 16 6644 26
rect 6896 16 6960 26
rect 7212 16 7276 26
rect 7528 16 7592 26
rect 7844 16 7908 26
rect 8160 16 8224 26
rect 8476 16 8540 26
rect 8792 16 8856 26
rect 9108 16 9172 26
rect 9424 16 9488 26
rect 9740 16 9804 26
rect 10056 16 10120 26
rect 10372 16 10436 26
rect 10688 16 10752 26
rect 11004 16 11068 26
rect 11320 16 11384 26
rect 11636 16 11700 26
rect 11952 16 12016 26
rect 12268 16 12332 26
rect 12584 16 12648 26
rect 260 -18 274 16
rect 274 -18 310 16
rect 310 -18 324 16
rect 576 -18 590 16
rect 590 -18 626 16
rect 626 -18 640 16
rect 892 -18 906 16
rect 906 -18 942 16
rect 942 -18 956 16
rect 1208 -18 1222 16
rect 1222 -18 1258 16
rect 1258 -18 1272 16
rect 1524 -18 1538 16
rect 1538 -18 1574 16
rect 1574 -18 1588 16
rect 1840 -18 1854 16
rect 1854 -18 1890 16
rect 1890 -18 1904 16
rect 2156 -18 2170 16
rect 2170 -18 2206 16
rect 2206 -18 2220 16
rect 2472 -18 2486 16
rect 2486 -18 2522 16
rect 2522 -18 2536 16
rect 2788 -18 2802 16
rect 2802 -18 2838 16
rect 2838 -18 2852 16
rect 3104 -18 3118 16
rect 3118 -18 3154 16
rect 3154 -18 3168 16
rect 3420 -18 3434 16
rect 3434 -18 3470 16
rect 3470 -18 3484 16
rect 3736 -18 3750 16
rect 3750 -18 3786 16
rect 3786 -18 3800 16
rect 4052 -18 4066 16
rect 4066 -18 4102 16
rect 4102 -18 4116 16
rect 4368 -18 4382 16
rect 4382 -18 4418 16
rect 4418 -18 4432 16
rect 4684 -18 4698 16
rect 4698 -18 4734 16
rect 4734 -18 4748 16
rect 5000 -18 5014 16
rect 5014 -18 5050 16
rect 5050 -18 5064 16
rect 5316 -18 5330 16
rect 5330 -18 5366 16
rect 5366 -18 5380 16
rect 5632 -18 5646 16
rect 5646 -18 5682 16
rect 5682 -18 5696 16
rect 5948 -18 5962 16
rect 5962 -18 5998 16
rect 5998 -18 6012 16
rect 6264 -18 6278 16
rect 6278 -18 6314 16
rect 6314 -18 6328 16
rect 6580 -18 6594 16
rect 6594 -18 6630 16
rect 6630 -18 6644 16
rect 6896 -18 6910 16
rect 6910 -18 6946 16
rect 6946 -18 6960 16
rect 7212 -18 7226 16
rect 7226 -18 7262 16
rect 7262 -18 7276 16
rect 7528 -18 7542 16
rect 7542 -18 7578 16
rect 7578 -18 7592 16
rect 7844 -18 7858 16
rect 7858 -18 7894 16
rect 7894 -18 7908 16
rect 8160 -18 8174 16
rect 8174 -18 8210 16
rect 8210 -18 8224 16
rect 8476 -18 8490 16
rect 8490 -18 8526 16
rect 8526 -18 8540 16
rect 8792 -18 8806 16
rect 8806 -18 8842 16
rect 8842 -18 8856 16
rect 9108 -18 9122 16
rect 9122 -18 9158 16
rect 9158 -18 9172 16
rect 9424 -18 9438 16
rect 9438 -18 9474 16
rect 9474 -18 9488 16
rect 9740 -18 9754 16
rect 9754 -18 9790 16
rect 9790 -18 9804 16
rect 10056 -18 10070 16
rect 10070 -18 10106 16
rect 10106 -18 10120 16
rect 10372 -18 10386 16
rect 10386 -18 10422 16
rect 10422 -18 10436 16
rect 10688 -18 10702 16
rect 10702 -18 10738 16
rect 10738 -18 10752 16
rect 11004 -18 11018 16
rect 11018 -18 11054 16
rect 11054 -18 11068 16
rect 11320 -18 11334 16
rect 11334 -18 11370 16
rect 11370 -18 11384 16
rect 11636 -18 11650 16
rect 11650 -18 11686 16
rect 11686 -18 11700 16
rect 11952 -18 11966 16
rect 11966 -18 12002 16
rect 12002 -18 12016 16
rect 12268 -18 12282 16
rect 12282 -18 12318 16
rect 12318 -18 12332 16
rect 12584 -18 12598 16
rect 12598 -18 12634 16
rect 12634 -18 12648 16
rect 260 -28 324 -18
rect 576 -28 640 -18
rect 892 -28 956 -18
rect 1208 -28 1272 -18
rect 1524 -28 1588 -18
rect 1840 -28 1904 -18
rect 2156 -28 2220 -18
rect 2472 -28 2536 -18
rect 2788 -28 2852 -18
rect 3104 -28 3168 -18
rect 3420 -28 3484 -18
rect 3736 -28 3800 -18
rect 4052 -28 4116 -18
rect 4368 -28 4432 -18
rect 4684 -28 4748 -18
rect 5000 -28 5064 -18
rect 5316 -28 5380 -18
rect 5632 -28 5696 -18
rect 5948 -28 6012 -18
rect 6264 -28 6328 -18
rect 6580 -28 6644 -18
rect 6896 -28 6960 -18
rect 7212 -28 7276 -18
rect 7528 -28 7592 -18
rect 7844 -28 7908 -18
rect 8160 -28 8224 -18
rect 8476 -28 8540 -18
rect 8792 -28 8856 -18
rect 9108 -28 9172 -18
rect 9424 -28 9488 -18
rect 9740 -28 9804 -18
rect 10056 -28 10120 -18
rect 10372 -28 10436 -18
rect 10688 -28 10752 -18
rect 11004 -28 11068 -18
rect 11320 -28 11384 -18
rect 11636 -28 11700 -18
rect 11952 -28 12016 -18
rect 12268 -28 12332 -18
rect 12584 -28 12648 -18
<< metal2 >>
rect 110 4632 158 4890
rect 268 4858 316 4890
rect 254 4852 330 4858
rect 254 4798 260 4852
rect 324 4798 330 4852
rect 254 4792 330 4798
rect 268 4632 316 4792
rect 426 4632 474 4890
rect 584 4858 632 4890
rect 570 4852 646 4858
rect 570 4798 576 4852
rect 640 4798 646 4852
rect 570 4792 646 4798
rect 584 4632 632 4792
rect 742 4632 790 4890
rect 900 4858 948 4890
rect 886 4852 962 4858
rect 886 4798 892 4852
rect 956 4798 962 4852
rect 886 4792 962 4798
rect 900 4632 948 4792
rect 1058 4632 1106 4890
rect 1216 4858 1264 4890
rect 1202 4852 1278 4858
rect 1202 4798 1208 4852
rect 1272 4798 1278 4852
rect 1202 4792 1278 4798
rect 1216 4632 1264 4792
rect 1374 4632 1422 4890
rect 1532 4858 1580 4890
rect 1518 4852 1594 4858
rect 1518 4798 1524 4852
rect 1588 4798 1594 4852
rect 1518 4792 1594 4798
rect 1532 4632 1580 4792
rect 1690 4632 1738 4890
rect 1848 4858 1896 4890
rect 1834 4852 1910 4858
rect 1834 4798 1840 4852
rect 1904 4798 1910 4852
rect 1834 4792 1910 4798
rect 1848 4632 1896 4792
rect 2006 4632 2054 4890
rect 2164 4858 2212 4890
rect 2150 4852 2226 4858
rect 2150 4798 2156 4852
rect 2220 4798 2226 4852
rect 2150 4792 2226 4798
rect 2164 4632 2212 4792
rect 2322 4632 2370 4890
rect 2480 4858 2528 4890
rect 2466 4852 2542 4858
rect 2466 4798 2472 4852
rect 2536 4798 2542 4852
rect 2466 4792 2542 4798
rect 2480 4632 2528 4792
rect 2638 4632 2686 4890
rect 2796 4858 2844 4890
rect 2782 4852 2858 4858
rect 2782 4798 2788 4852
rect 2852 4798 2858 4852
rect 2782 4792 2858 4798
rect 2796 4632 2844 4792
rect 2954 4632 3002 4890
rect 3112 4858 3160 4890
rect 3098 4852 3174 4858
rect 3098 4798 3104 4852
rect 3168 4798 3174 4852
rect 3098 4792 3174 4798
rect 3112 4632 3160 4792
rect 3270 4632 3318 4890
rect 3428 4858 3476 4890
rect 3414 4852 3490 4858
rect 3414 4798 3420 4852
rect 3484 4798 3490 4852
rect 3414 4792 3490 4798
rect 3428 4632 3476 4792
rect 3586 4632 3634 4890
rect 3744 4858 3792 4890
rect 3730 4852 3806 4858
rect 3730 4798 3736 4852
rect 3800 4798 3806 4852
rect 3730 4792 3806 4798
rect 3744 4632 3792 4792
rect 3902 4632 3950 4890
rect 4060 4858 4108 4890
rect 4046 4852 4122 4858
rect 4046 4798 4052 4852
rect 4116 4798 4122 4852
rect 4046 4792 4122 4798
rect 4060 4632 4108 4792
rect 4218 4632 4266 4890
rect 4376 4858 4424 4890
rect 4362 4852 4438 4858
rect 4362 4798 4368 4852
rect 4432 4798 4438 4852
rect 4362 4792 4438 4798
rect 4376 4632 4424 4792
rect 4534 4632 4582 4890
rect 4692 4858 4740 4890
rect 4678 4852 4754 4858
rect 4678 4798 4684 4852
rect 4748 4798 4754 4852
rect 4678 4792 4754 4798
rect 4692 4632 4740 4792
rect 4850 4632 4898 4890
rect 5008 4858 5056 4890
rect 4994 4852 5070 4858
rect 4994 4798 5000 4852
rect 5064 4798 5070 4852
rect 4994 4792 5070 4798
rect 5008 4632 5056 4792
rect 5166 4632 5214 4890
rect 5324 4858 5372 4890
rect 5310 4852 5386 4858
rect 5310 4798 5316 4852
rect 5380 4798 5386 4852
rect 5310 4792 5386 4798
rect 5324 4632 5372 4792
rect 5482 4632 5530 4890
rect 5640 4858 5688 4890
rect 5626 4852 5702 4858
rect 5626 4798 5632 4852
rect 5696 4798 5702 4852
rect 5626 4792 5702 4798
rect 5640 4632 5688 4792
rect 5798 4632 5846 4890
rect 5956 4858 6004 4890
rect 5942 4852 6018 4858
rect 5942 4798 5948 4852
rect 6012 4798 6018 4852
rect 5942 4792 6018 4798
rect 5956 4632 6004 4792
rect 6114 4632 6162 4890
rect 6272 4858 6320 4890
rect 6258 4852 6334 4858
rect 6258 4798 6264 4852
rect 6328 4798 6334 4852
rect 6258 4792 6334 4798
rect 6272 4632 6320 4792
rect 6430 4632 6478 4890
rect 6588 4858 6636 4890
rect 6574 4852 6650 4858
rect 6574 4798 6580 4852
rect 6644 4798 6650 4852
rect 6574 4792 6650 4798
rect 6588 4632 6636 4792
rect 6746 4632 6794 4890
rect 6904 4858 6952 4890
rect 6890 4852 6966 4858
rect 6890 4798 6896 4852
rect 6960 4798 6966 4852
rect 6890 4792 6966 4798
rect 6904 4632 6952 4792
rect 7062 4632 7110 4890
rect 7220 4858 7268 4890
rect 7206 4852 7282 4858
rect 7206 4798 7212 4852
rect 7276 4798 7282 4852
rect 7206 4792 7282 4798
rect 7220 4632 7268 4792
rect 7378 4632 7426 4890
rect 7536 4858 7584 4890
rect 7522 4852 7598 4858
rect 7522 4798 7528 4852
rect 7592 4798 7598 4852
rect 7522 4792 7598 4798
rect 7536 4632 7584 4792
rect 7694 4632 7742 4890
rect 7852 4858 7900 4890
rect 7838 4852 7914 4858
rect 7838 4798 7844 4852
rect 7908 4798 7914 4852
rect 7838 4792 7914 4798
rect 7852 4632 7900 4792
rect 8010 4632 8058 4890
rect 8168 4858 8216 4890
rect 8154 4852 8230 4858
rect 8154 4798 8160 4852
rect 8224 4798 8230 4852
rect 8154 4792 8230 4798
rect 8168 4632 8216 4792
rect 8326 4632 8374 4890
rect 8484 4858 8532 4890
rect 8470 4852 8546 4858
rect 8470 4798 8476 4852
rect 8540 4798 8546 4852
rect 8470 4792 8546 4798
rect 8484 4632 8532 4792
rect 8642 4632 8690 4890
rect 8800 4858 8848 4890
rect 8786 4852 8862 4858
rect 8786 4798 8792 4852
rect 8856 4798 8862 4852
rect 8786 4792 8862 4798
rect 8800 4632 8848 4792
rect 8958 4632 9006 4890
rect 9116 4858 9164 4890
rect 9102 4852 9178 4858
rect 9102 4798 9108 4852
rect 9172 4798 9178 4852
rect 9102 4792 9178 4798
rect 9116 4632 9164 4792
rect 9274 4632 9322 4890
rect 9432 4858 9480 4890
rect 9418 4852 9494 4858
rect 9418 4798 9424 4852
rect 9488 4798 9494 4852
rect 9418 4792 9494 4798
rect 9432 4632 9480 4792
rect 9590 4632 9638 4890
rect 9748 4858 9796 4890
rect 9734 4852 9810 4858
rect 9734 4798 9740 4852
rect 9804 4798 9810 4852
rect 9734 4792 9810 4798
rect 9748 4632 9796 4792
rect 9906 4632 9954 4890
rect 10064 4858 10112 4890
rect 10050 4852 10126 4858
rect 10050 4798 10056 4852
rect 10120 4798 10126 4852
rect 10050 4792 10126 4798
rect 10064 4632 10112 4792
rect 10222 4632 10270 4890
rect 10380 4858 10428 4890
rect 10366 4852 10442 4858
rect 10366 4798 10372 4852
rect 10436 4798 10442 4852
rect 10366 4792 10442 4798
rect 10380 4632 10428 4792
rect 10538 4632 10586 4890
rect 10696 4858 10744 4890
rect 10682 4852 10758 4858
rect 10682 4798 10688 4852
rect 10752 4798 10758 4852
rect 10682 4792 10758 4798
rect 10696 4632 10744 4792
rect 10854 4632 10902 4890
rect 11012 4858 11060 4890
rect 10998 4852 11074 4858
rect 10998 4798 11004 4852
rect 11068 4798 11074 4852
rect 10998 4792 11074 4798
rect 11012 4632 11060 4792
rect 11170 4632 11218 4890
rect 11328 4858 11376 4890
rect 11314 4852 11390 4858
rect 11314 4798 11320 4852
rect 11384 4798 11390 4852
rect 11314 4792 11390 4798
rect 11328 4632 11376 4792
rect 11486 4632 11534 4890
rect 11644 4858 11692 4890
rect 11630 4852 11706 4858
rect 11630 4798 11636 4852
rect 11700 4798 11706 4852
rect 11630 4792 11706 4798
rect 11644 4632 11692 4792
rect 11802 4632 11850 4890
rect 11960 4858 12008 4890
rect 11946 4852 12022 4858
rect 11946 4798 11952 4852
rect 12016 4798 12022 4852
rect 11946 4792 12022 4798
rect 11960 4632 12008 4792
rect 12118 4632 12166 4890
rect 12276 4858 12324 4890
rect 12262 4852 12338 4858
rect 12262 4798 12268 4852
rect 12332 4798 12338 4852
rect 12262 4792 12338 4798
rect 12276 4632 12324 4792
rect 12434 4632 12482 4890
rect 12592 4858 12640 4890
rect 12578 4852 12654 4858
rect 12578 4798 12584 4852
rect 12648 4798 12654 4852
rect 12578 4792 12654 4798
rect 12592 4632 12640 4792
rect 12750 4750 12798 4890
rect 12744 4632 12798 4750
rect 98 4622 172 4632
rect 98 3844 108 4622
rect 164 3844 172 4622
rect 98 3834 172 3844
rect 256 4622 328 4632
rect 256 3840 266 4622
rect 322 3840 328 4622
rect 110 3722 158 3834
rect 256 3830 328 3840
rect 412 4622 488 4632
rect 412 3840 422 4622
rect 478 3840 488 4622
rect 412 3830 488 3840
rect 572 4622 644 4632
rect 572 3840 582 4622
rect 638 3840 644 4622
rect 572 3830 644 3840
rect 728 4622 804 4632
rect 728 3840 738 4622
rect 794 3840 804 4622
rect 728 3830 804 3840
rect 888 4622 960 4632
rect 888 3840 898 4622
rect 954 3840 960 4622
rect 888 3830 960 3840
rect 1044 4622 1120 4632
rect 1044 3840 1054 4622
rect 1110 3840 1120 4622
rect 1044 3830 1120 3840
rect 1204 4622 1276 4632
rect 1204 3840 1214 4622
rect 1270 3840 1276 4622
rect 1204 3830 1276 3840
rect 1360 4622 1436 4632
rect 1360 3840 1370 4622
rect 1426 3840 1436 4622
rect 1360 3830 1436 3840
rect 1520 4622 1592 4632
rect 1520 3840 1530 4622
rect 1586 3840 1592 4622
rect 1520 3830 1592 3840
rect 1676 4622 1752 4632
rect 1676 3840 1686 4622
rect 1742 3840 1752 4622
rect 1676 3830 1752 3840
rect 1836 4622 1908 4632
rect 1836 3840 1846 4622
rect 1902 3840 1908 4622
rect 1836 3830 1908 3840
rect 1992 4622 2068 4632
rect 1992 3840 2002 4622
rect 2058 3840 2068 4622
rect 1992 3830 2068 3840
rect 2152 4622 2224 4632
rect 2152 3840 2162 4622
rect 2218 3840 2224 4622
rect 2152 3830 2224 3840
rect 2308 4622 2384 4632
rect 2308 3840 2318 4622
rect 2374 3840 2384 4622
rect 2308 3830 2384 3840
rect 2468 4622 2540 4632
rect 2468 3840 2478 4622
rect 2534 3840 2540 4622
rect 2468 3830 2540 3840
rect 2624 4622 2700 4632
rect 2624 3840 2634 4622
rect 2690 3840 2700 4622
rect 2624 3830 2700 3840
rect 2784 4622 2856 4632
rect 2784 3840 2794 4622
rect 2850 3840 2856 4622
rect 2784 3830 2856 3840
rect 2940 4622 3016 4632
rect 2940 3840 2950 4622
rect 3006 3840 3016 4622
rect 2940 3830 3016 3840
rect 3100 4622 3172 4632
rect 3100 3840 3110 4622
rect 3166 3840 3172 4622
rect 3100 3830 3172 3840
rect 3256 4622 3332 4632
rect 3256 3840 3266 4622
rect 3322 3840 3332 4622
rect 3256 3830 3332 3840
rect 3416 4622 3488 4632
rect 3416 3840 3426 4622
rect 3482 3840 3488 4622
rect 3416 3830 3488 3840
rect 3572 4622 3648 4632
rect 3572 3840 3582 4622
rect 3638 3840 3648 4622
rect 3572 3830 3648 3840
rect 3732 4622 3804 4632
rect 3732 3840 3742 4622
rect 3798 3840 3804 4622
rect 3732 3830 3804 3840
rect 3888 4622 3964 4632
rect 3888 3840 3898 4622
rect 3954 3840 3964 4622
rect 3888 3830 3964 3840
rect 4048 4622 4120 4632
rect 4048 3840 4058 4622
rect 4114 3840 4120 4622
rect 4048 3830 4120 3840
rect 4204 4622 4280 4632
rect 4204 3840 4214 4622
rect 4270 3840 4280 4622
rect 4204 3830 4280 3840
rect 4364 4622 4436 4632
rect 4364 3840 4374 4622
rect 4430 3840 4436 4622
rect 4364 3830 4436 3840
rect 4520 4622 4596 4632
rect 4520 3840 4530 4622
rect 4586 3840 4596 4622
rect 4520 3830 4596 3840
rect 4680 4622 4752 4632
rect 4680 3840 4690 4622
rect 4746 3840 4752 4622
rect 4680 3830 4752 3840
rect 4836 4622 4912 4632
rect 4836 3840 4846 4622
rect 4902 3840 4912 4622
rect 4836 3830 4912 3840
rect 4996 4622 5068 4632
rect 4996 3840 5006 4622
rect 5062 3840 5068 4622
rect 4996 3830 5068 3840
rect 5152 4622 5228 4632
rect 5152 3840 5162 4622
rect 5218 3840 5228 4622
rect 5152 3830 5228 3840
rect 5312 4622 5384 4632
rect 5312 3840 5322 4622
rect 5378 3840 5384 4622
rect 5312 3830 5384 3840
rect 5468 4622 5544 4632
rect 5468 3840 5478 4622
rect 5534 3840 5544 4622
rect 5468 3830 5544 3840
rect 5628 4622 5700 4632
rect 5628 3840 5638 4622
rect 5694 3840 5700 4622
rect 5628 3830 5700 3840
rect 5784 4622 5860 4632
rect 5784 3840 5794 4622
rect 5850 3840 5860 4622
rect 5784 3830 5860 3840
rect 5944 4622 6016 4632
rect 5944 3840 5954 4622
rect 6010 3840 6016 4622
rect 5944 3830 6016 3840
rect 6100 4622 6176 4632
rect 6100 3840 6110 4622
rect 6166 3840 6176 4622
rect 6100 3830 6176 3840
rect 6260 4622 6332 4632
rect 6260 3840 6270 4622
rect 6326 3840 6332 4622
rect 6260 3830 6332 3840
rect 6416 4622 6492 4632
rect 6416 3840 6426 4622
rect 6482 3840 6492 4622
rect 6416 3830 6492 3840
rect 6576 4622 6648 4632
rect 6576 3840 6586 4622
rect 6642 3840 6648 4622
rect 6576 3830 6648 3840
rect 6732 4622 6808 4632
rect 6732 3840 6742 4622
rect 6798 3840 6808 4622
rect 6732 3830 6808 3840
rect 6892 4622 6964 4632
rect 6892 3840 6902 4622
rect 6958 3840 6964 4622
rect 6892 3830 6964 3840
rect 7048 4622 7124 4632
rect 7048 3840 7058 4622
rect 7114 3840 7124 4622
rect 7048 3830 7124 3840
rect 7208 4622 7280 4632
rect 7208 3840 7218 4622
rect 7274 3840 7280 4622
rect 7208 3830 7280 3840
rect 7364 4622 7440 4632
rect 7364 3840 7374 4622
rect 7430 3840 7440 4622
rect 7364 3830 7440 3840
rect 7524 4622 7596 4632
rect 7524 3840 7534 4622
rect 7590 3840 7596 4622
rect 7524 3830 7596 3840
rect 7680 4622 7756 4632
rect 7680 3840 7690 4622
rect 7746 3840 7756 4622
rect 7680 3830 7756 3840
rect 7840 4622 7912 4632
rect 7840 3840 7850 4622
rect 7906 3840 7912 4622
rect 7840 3830 7912 3840
rect 7996 4622 8072 4632
rect 7996 3840 8006 4622
rect 8062 3840 8072 4622
rect 7996 3830 8072 3840
rect 8156 4622 8228 4632
rect 8156 3840 8166 4622
rect 8222 3840 8228 4622
rect 8156 3830 8228 3840
rect 8312 4622 8388 4632
rect 8312 3840 8322 4622
rect 8378 3840 8388 4622
rect 8312 3830 8388 3840
rect 8472 4622 8544 4632
rect 8472 3840 8482 4622
rect 8538 3840 8544 4622
rect 8472 3830 8544 3840
rect 8628 4622 8704 4632
rect 8628 3840 8638 4622
rect 8694 3840 8704 4622
rect 8628 3830 8704 3840
rect 8788 4622 8860 4632
rect 8788 3840 8798 4622
rect 8854 3840 8860 4622
rect 8788 3830 8860 3840
rect 8944 4622 9020 4632
rect 8944 3840 8954 4622
rect 9010 3840 9020 4622
rect 8944 3830 9020 3840
rect 9104 4622 9176 4632
rect 9104 3840 9114 4622
rect 9170 3840 9176 4622
rect 9104 3830 9176 3840
rect 9260 4622 9336 4632
rect 9260 3840 9270 4622
rect 9326 3840 9336 4622
rect 9260 3830 9336 3840
rect 9420 4622 9492 4632
rect 9420 3840 9430 4622
rect 9486 3840 9492 4622
rect 9420 3830 9492 3840
rect 9576 4622 9652 4632
rect 9576 3840 9586 4622
rect 9642 3840 9652 4622
rect 9576 3830 9652 3840
rect 9736 4622 9808 4632
rect 9736 3840 9746 4622
rect 9802 3840 9808 4622
rect 9736 3830 9808 3840
rect 9892 4622 9968 4632
rect 9892 3840 9902 4622
rect 9958 3840 9968 4622
rect 9892 3830 9968 3840
rect 10052 4622 10124 4632
rect 10052 3840 10062 4622
rect 10118 3840 10124 4622
rect 10052 3830 10124 3840
rect 10208 4622 10284 4632
rect 10208 3840 10218 4622
rect 10274 3840 10284 4622
rect 10208 3830 10284 3840
rect 10368 4622 10440 4632
rect 10368 3840 10378 4622
rect 10434 3840 10440 4622
rect 10368 3830 10440 3840
rect 10524 4622 10600 4632
rect 10524 3840 10534 4622
rect 10590 3840 10600 4622
rect 10524 3830 10600 3840
rect 10684 4622 10756 4632
rect 10684 3840 10694 4622
rect 10750 3840 10756 4622
rect 10684 3830 10756 3840
rect 10840 4622 10916 4632
rect 10840 3840 10850 4622
rect 10906 3840 10916 4622
rect 10840 3830 10916 3840
rect 11000 4622 11072 4632
rect 11000 3840 11010 4622
rect 11066 3840 11072 4622
rect 11000 3830 11072 3840
rect 11156 4622 11232 4632
rect 11156 3840 11166 4622
rect 11222 3840 11232 4622
rect 11156 3830 11232 3840
rect 11316 4622 11388 4632
rect 11316 3840 11326 4622
rect 11382 3840 11388 4622
rect 11316 3830 11388 3840
rect 11472 4622 11548 4632
rect 11472 3840 11482 4622
rect 11538 3840 11548 4622
rect 11472 3830 11548 3840
rect 11632 4622 11704 4632
rect 11632 3840 11642 4622
rect 11698 3840 11704 4622
rect 11632 3830 11704 3840
rect 11788 4622 11864 4632
rect 11788 3840 11798 4622
rect 11854 3840 11864 4622
rect 11788 3830 11864 3840
rect 11948 4622 12020 4632
rect 11948 3840 11958 4622
rect 12014 3840 12020 4622
rect 11948 3830 12020 3840
rect 12104 4622 12180 4632
rect 12104 3840 12114 4622
rect 12170 3840 12180 4622
rect 12104 3830 12180 3840
rect 12264 4622 12336 4632
rect 12264 3840 12274 4622
rect 12330 3840 12336 4622
rect 12264 3830 12336 3840
rect 12420 4622 12496 4632
rect 12420 3840 12430 4622
rect 12486 3840 12496 4622
rect 12420 3830 12496 3840
rect 12580 4622 12652 4632
rect 12580 3840 12590 4622
rect 12646 3840 12652 4622
rect 12580 3830 12652 3840
rect 12736 4622 12812 4632
rect 12736 3844 12744 4622
rect 12736 3840 12746 3844
rect 12802 3840 12812 4622
rect 12736 3830 12812 3840
rect 268 3722 316 3830
rect 426 3722 474 3830
rect 584 3722 632 3830
rect 742 3722 790 3830
rect 900 3722 948 3830
rect 1058 3722 1106 3830
rect 1216 3722 1264 3830
rect 1374 3722 1422 3830
rect 1532 3722 1580 3830
rect 1690 3722 1738 3830
rect 1848 3722 1896 3830
rect 2006 3722 2054 3830
rect 2164 3722 2212 3830
rect 2322 3722 2370 3830
rect 2480 3722 2528 3830
rect 2638 3722 2686 3830
rect 2796 3722 2844 3830
rect 2954 3722 3002 3830
rect 3112 3722 3160 3830
rect 3270 3722 3318 3830
rect 3428 3722 3476 3830
rect 3586 3722 3634 3830
rect 3744 3722 3792 3830
rect 3902 3722 3950 3830
rect 4060 3722 4108 3830
rect 4218 3722 4266 3830
rect 4376 3722 4424 3830
rect 4534 3722 4582 3830
rect 4692 3722 4740 3830
rect 4850 3722 4898 3830
rect 5008 3722 5056 3830
rect 5166 3722 5214 3830
rect 5324 3722 5372 3830
rect 5482 3722 5530 3830
rect 5640 3722 5688 3830
rect 5798 3722 5846 3830
rect 5956 3722 6004 3830
rect 6114 3722 6162 3830
rect 6272 3722 6320 3830
rect 6430 3722 6478 3830
rect 6588 3722 6636 3830
rect 6746 3722 6794 3830
rect 6904 3722 6952 3830
rect 7062 3722 7110 3830
rect 7220 3722 7268 3830
rect 7378 3722 7426 3830
rect 7536 3722 7584 3830
rect 7694 3722 7742 3830
rect 7852 3722 7900 3830
rect 8010 3722 8058 3830
rect 8168 3722 8216 3830
rect 8326 3722 8374 3830
rect 8484 3722 8532 3830
rect 8642 3722 8690 3830
rect 8800 3722 8848 3830
rect 8958 3722 9006 3830
rect 9116 3722 9164 3830
rect 9274 3722 9322 3830
rect 9432 3722 9480 3830
rect 9590 3722 9638 3830
rect 9748 3722 9796 3830
rect 9906 3722 9954 3830
rect 10064 3722 10112 3830
rect 10222 3722 10270 3830
rect 10380 3722 10428 3830
rect 10538 3722 10586 3830
rect 10696 3722 10744 3830
rect 10854 3722 10902 3830
rect 11012 3722 11060 3830
rect 11170 3722 11218 3830
rect 11328 3722 11376 3830
rect 11486 3722 11534 3830
rect 11644 3722 11692 3830
rect 11802 3722 11850 3830
rect 11960 3722 12008 3830
rect 12118 3722 12166 3830
rect 12276 3722 12324 3830
rect 12434 3722 12482 3830
rect 12592 3722 12640 3830
rect 12744 3722 12798 3830
rect 98 3714 172 3722
rect 98 3712 110 3714
rect 162 3712 172 3714
rect 98 2934 108 3712
rect 164 2934 172 3712
rect 98 2932 110 2934
rect 162 2932 172 2934
rect 98 2924 172 2932
rect 256 3712 328 3722
rect 256 2930 266 3712
rect 322 2930 328 3712
rect 110 2812 158 2924
rect 256 2920 328 2930
rect 412 3714 488 3722
rect 412 3712 426 3714
rect 412 2930 422 3712
rect 478 2930 488 3714
rect 412 2920 488 2930
rect 572 3712 644 3722
rect 572 2930 582 3712
rect 638 2930 644 3712
rect 572 2920 644 2930
rect 728 3714 804 3722
rect 728 3712 742 3714
rect 728 2930 738 3712
rect 794 2930 804 3714
rect 728 2920 804 2930
rect 888 3712 960 3722
rect 888 2930 898 3712
rect 954 2930 960 3712
rect 888 2920 960 2930
rect 1044 3714 1120 3722
rect 1044 3712 1058 3714
rect 1044 2930 1054 3712
rect 1110 2930 1120 3714
rect 1044 2920 1120 2930
rect 1204 3712 1276 3722
rect 1204 2930 1214 3712
rect 1270 2930 1276 3712
rect 1204 2920 1276 2930
rect 1360 3714 1436 3722
rect 1360 3712 1374 3714
rect 1360 2930 1370 3712
rect 1426 2930 1436 3714
rect 1360 2920 1436 2930
rect 1520 3712 1592 3722
rect 1520 2930 1530 3712
rect 1586 2930 1592 3712
rect 1520 2920 1592 2930
rect 1676 3714 1752 3722
rect 1676 3712 1690 3714
rect 1676 2930 1686 3712
rect 1742 2930 1752 3714
rect 1676 2920 1752 2930
rect 1836 3712 1908 3722
rect 1836 2930 1846 3712
rect 1902 2930 1908 3712
rect 1836 2920 1908 2930
rect 1992 3714 2068 3722
rect 1992 3712 2006 3714
rect 1992 2930 2002 3712
rect 2058 2930 2068 3714
rect 1992 2920 2068 2930
rect 2152 3712 2224 3722
rect 2152 2930 2162 3712
rect 2218 2930 2224 3712
rect 2152 2920 2224 2930
rect 2308 3714 2384 3722
rect 2308 3712 2322 3714
rect 2308 2930 2318 3712
rect 2374 2930 2384 3714
rect 2308 2920 2384 2930
rect 2468 3712 2540 3722
rect 2468 2930 2478 3712
rect 2534 2930 2540 3712
rect 2468 2920 2540 2930
rect 2624 3714 2700 3722
rect 2624 3712 2638 3714
rect 2624 2930 2634 3712
rect 2690 2930 2700 3714
rect 2624 2920 2700 2930
rect 2784 3712 2856 3722
rect 2784 2930 2794 3712
rect 2850 2930 2856 3712
rect 2784 2920 2856 2930
rect 2940 3714 3016 3722
rect 2940 3712 2954 3714
rect 2940 2930 2950 3712
rect 3006 2930 3016 3714
rect 2940 2920 3016 2930
rect 3100 3712 3172 3722
rect 3100 2930 3110 3712
rect 3166 2930 3172 3712
rect 3100 2920 3172 2930
rect 3256 3714 3332 3722
rect 3256 3712 3270 3714
rect 3256 2930 3266 3712
rect 3322 2930 3332 3714
rect 3256 2920 3332 2930
rect 3416 3712 3488 3722
rect 3416 2930 3426 3712
rect 3482 2930 3488 3712
rect 3416 2920 3488 2930
rect 3572 3714 3648 3722
rect 3572 3712 3586 3714
rect 3572 2930 3582 3712
rect 3638 2930 3648 3714
rect 3572 2920 3648 2930
rect 3732 3712 3804 3722
rect 3732 2930 3742 3712
rect 3798 2930 3804 3712
rect 3732 2920 3804 2930
rect 3888 3714 3964 3722
rect 3888 3712 3902 3714
rect 3888 2930 3898 3712
rect 3954 2930 3964 3714
rect 3888 2920 3964 2930
rect 4048 3712 4120 3722
rect 4048 2930 4058 3712
rect 4114 2930 4120 3712
rect 4048 2920 4120 2930
rect 4204 3714 4280 3722
rect 4204 3712 4218 3714
rect 4204 2930 4214 3712
rect 4270 2930 4280 3714
rect 4204 2920 4280 2930
rect 4364 3712 4436 3722
rect 4364 2930 4374 3712
rect 4430 2930 4436 3712
rect 4364 2920 4436 2930
rect 4520 3714 4596 3722
rect 4520 3712 4534 3714
rect 4520 2930 4530 3712
rect 4586 2930 4596 3714
rect 4520 2920 4596 2930
rect 4680 3712 4752 3722
rect 4680 2930 4690 3712
rect 4746 2930 4752 3712
rect 4680 2920 4752 2930
rect 4836 3714 4912 3722
rect 4836 3712 4850 3714
rect 4836 2930 4846 3712
rect 4902 2930 4912 3714
rect 4836 2920 4912 2930
rect 4996 3712 5068 3722
rect 4996 2930 5006 3712
rect 5062 2930 5068 3712
rect 4996 2920 5068 2930
rect 5152 3714 5228 3722
rect 5152 3712 5166 3714
rect 5152 2930 5162 3712
rect 5218 2930 5228 3714
rect 5152 2920 5228 2930
rect 5312 3712 5384 3722
rect 5312 2930 5322 3712
rect 5378 2930 5384 3712
rect 5312 2920 5384 2930
rect 5468 3714 5544 3722
rect 5468 3712 5482 3714
rect 5468 2930 5478 3712
rect 5534 2930 5544 3714
rect 5468 2920 5544 2930
rect 5628 3712 5700 3722
rect 5628 2930 5638 3712
rect 5694 2930 5700 3712
rect 5628 2920 5700 2930
rect 5784 3714 5860 3722
rect 5784 3712 5798 3714
rect 5784 2930 5794 3712
rect 5850 2930 5860 3714
rect 5784 2920 5860 2930
rect 5944 3712 6016 3722
rect 5944 2930 5954 3712
rect 6010 2930 6016 3712
rect 5944 2920 6016 2930
rect 6100 3714 6176 3722
rect 6100 3712 6114 3714
rect 6100 2930 6110 3712
rect 6166 2930 6176 3714
rect 6100 2920 6176 2930
rect 6260 3712 6332 3722
rect 6260 2930 6270 3712
rect 6326 2930 6332 3712
rect 6260 2920 6332 2930
rect 6416 3714 6492 3722
rect 6416 3712 6430 3714
rect 6416 2930 6426 3712
rect 6482 2930 6492 3714
rect 6416 2920 6492 2930
rect 6576 3712 6648 3722
rect 6576 2930 6586 3712
rect 6642 2930 6648 3712
rect 6576 2920 6648 2930
rect 6732 3714 6808 3722
rect 6732 3712 6746 3714
rect 6732 2930 6742 3712
rect 6798 2930 6808 3714
rect 6732 2920 6808 2930
rect 6892 3712 6964 3722
rect 6892 2930 6902 3712
rect 6958 2930 6964 3712
rect 6892 2920 6964 2930
rect 7048 3714 7124 3722
rect 7048 3712 7062 3714
rect 7048 2930 7058 3712
rect 7114 2930 7124 3714
rect 7048 2920 7124 2930
rect 7208 3712 7280 3722
rect 7208 2930 7218 3712
rect 7274 2930 7280 3712
rect 7208 2920 7280 2930
rect 7364 3714 7440 3722
rect 7364 3712 7378 3714
rect 7364 2930 7374 3712
rect 7430 2930 7440 3714
rect 7364 2920 7440 2930
rect 7524 3712 7596 3722
rect 7524 2930 7534 3712
rect 7590 2930 7596 3712
rect 7524 2920 7596 2930
rect 7680 3714 7756 3722
rect 7680 3712 7694 3714
rect 7680 2930 7690 3712
rect 7746 2930 7756 3714
rect 7680 2920 7756 2930
rect 7840 3712 7912 3722
rect 7840 2930 7850 3712
rect 7906 2930 7912 3712
rect 7840 2920 7912 2930
rect 7996 3714 8072 3722
rect 7996 3712 8010 3714
rect 7996 2930 8006 3712
rect 8062 2930 8072 3714
rect 7996 2920 8072 2930
rect 8156 3712 8228 3722
rect 8156 2930 8166 3712
rect 8222 2930 8228 3712
rect 8156 2920 8228 2930
rect 8312 3714 8388 3722
rect 8312 3712 8326 3714
rect 8312 2930 8322 3712
rect 8378 2930 8388 3714
rect 8312 2920 8388 2930
rect 8472 3712 8544 3722
rect 8472 2930 8482 3712
rect 8538 2930 8544 3712
rect 8472 2920 8544 2930
rect 8628 3714 8704 3722
rect 8628 3712 8642 3714
rect 8628 2930 8638 3712
rect 8694 2930 8704 3714
rect 8628 2920 8704 2930
rect 8788 3712 8860 3722
rect 8788 2930 8798 3712
rect 8854 2930 8860 3712
rect 8788 2920 8860 2930
rect 8944 3714 9020 3722
rect 8944 3712 8958 3714
rect 8944 2930 8954 3712
rect 9010 2930 9020 3714
rect 8944 2920 9020 2930
rect 9104 3712 9176 3722
rect 9104 2930 9114 3712
rect 9170 2930 9176 3712
rect 9104 2920 9176 2930
rect 9260 3714 9336 3722
rect 9260 3712 9274 3714
rect 9260 2930 9270 3712
rect 9326 2930 9336 3714
rect 9260 2920 9336 2930
rect 9420 3712 9492 3722
rect 9420 2930 9430 3712
rect 9486 2930 9492 3712
rect 9420 2920 9492 2930
rect 9576 3714 9652 3722
rect 9576 3712 9590 3714
rect 9576 2930 9586 3712
rect 9642 2930 9652 3714
rect 9576 2920 9652 2930
rect 9736 3712 9808 3722
rect 9736 2930 9746 3712
rect 9802 2930 9808 3712
rect 9736 2920 9808 2930
rect 9892 3714 9968 3722
rect 9892 3712 9906 3714
rect 9892 2930 9902 3712
rect 9958 2930 9968 3714
rect 9892 2920 9968 2930
rect 10052 3712 10124 3722
rect 10052 2930 10062 3712
rect 10118 2930 10124 3712
rect 10052 2920 10124 2930
rect 10208 3714 10284 3722
rect 10208 3712 10222 3714
rect 10208 2930 10218 3712
rect 10274 2930 10284 3714
rect 10208 2920 10284 2930
rect 10368 3712 10440 3722
rect 10368 2930 10378 3712
rect 10434 2930 10440 3712
rect 10368 2920 10440 2930
rect 10524 3714 10600 3722
rect 10524 3712 10538 3714
rect 10524 2930 10534 3712
rect 10590 2930 10600 3714
rect 10524 2920 10600 2930
rect 10684 3712 10756 3722
rect 10684 2930 10694 3712
rect 10750 2930 10756 3712
rect 10684 2920 10756 2930
rect 10840 3714 10916 3722
rect 10840 3712 10854 3714
rect 10840 2930 10850 3712
rect 10906 2930 10916 3714
rect 10840 2920 10916 2930
rect 11000 3712 11072 3722
rect 11000 2930 11010 3712
rect 11066 2930 11072 3712
rect 11000 2920 11072 2930
rect 11156 3714 11232 3722
rect 11156 3712 11170 3714
rect 11156 2930 11166 3712
rect 11222 2930 11232 3714
rect 11156 2920 11232 2930
rect 11316 3712 11388 3722
rect 11316 2930 11326 3712
rect 11382 2930 11388 3712
rect 11316 2920 11388 2930
rect 11472 3714 11548 3722
rect 11472 3712 11486 3714
rect 11472 2930 11482 3712
rect 11538 2930 11548 3714
rect 11472 2920 11548 2930
rect 11632 3712 11704 3722
rect 11632 2930 11642 3712
rect 11698 2930 11704 3712
rect 11632 2920 11704 2930
rect 11788 3714 11864 3722
rect 11788 3712 11802 3714
rect 11788 2930 11798 3712
rect 11854 2930 11864 3714
rect 11788 2920 11864 2930
rect 11948 3712 12020 3722
rect 11948 2930 11958 3712
rect 12014 2930 12020 3712
rect 11948 2920 12020 2930
rect 12104 3714 12180 3722
rect 12104 3712 12118 3714
rect 12104 2930 12114 3712
rect 12170 2930 12180 3714
rect 12104 2920 12180 2930
rect 12264 3712 12336 3722
rect 12264 2930 12274 3712
rect 12330 2930 12336 3712
rect 12264 2920 12336 2930
rect 12420 3714 12496 3722
rect 12420 3712 12434 3714
rect 12420 2930 12430 3712
rect 12486 2930 12496 3714
rect 12420 2920 12496 2930
rect 12580 3712 12652 3722
rect 12580 2930 12590 3712
rect 12646 2930 12652 3712
rect 12580 2920 12652 2930
rect 12736 3714 12812 3722
rect 12736 2932 12744 3714
rect 12796 3712 12812 3714
rect 12736 2930 12746 2932
rect 12802 2930 12812 3712
rect 12736 2920 12812 2930
rect 268 2812 316 2920
rect 426 2812 474 2920
rect 584 2812 632 2920
rect 742 2812 790 2920
rect 900 2812 948 2920
rect 1058 2812 1106 2920
rect 1216 2812 1264 2920
rect 1374 2812 1422 2920
rect 1532 2812 1580 2920
rect 1690 2812 1738 2920
rect 1848 2812 1896 2920
rect 2006 2812 2054 2920
rect 2164 2812 2212 2920
rect 2322 2812 2370 2920
rect 2480 2812 2528 2920
rect 2638 2812 2686 2920
rect 2796 2812 2844 2920
rect 2954 2812 3002 2920
rect 3112 2812 3160 2920
rect 3270 2812 3318 2920
rect 3428 2812 3476 2920
rect 3586 2812 3634 2920
rect 3744 2812 3792 2920
rect 3902 2812 3950 2920
rect 4060 2812 4108 2920
rect 4218 2812 4266 2920
rect 4376 2812 4424 2920
rect 4534 2812 4582 2920
rect 4692 2812 4740 2920
rect 4850 2812 4898 2920
rect 5008 2812 5056 2920
rect 5166 2812 5214 2920
rect 5324 2812 5372 2920
rect 5482 2812 5530 2920
rect 5640 2812 5688 2920
rect 5798 2812 5846 2920
rect 5956 2812 6004 2920
rect 6114 2812 6162 2920
rect 6272 2812 6320 2920
rect 6430 2812 6478 2920
rect 6588 2812 6636 2920
rect 6746 2812 6794 2920
rect 6904 2812 6952 2920
rect 7062 2812 7110 2920
rect 7220 2812 7268 2920
rect 7378 2812 7426 2920
rect 7536 2812 7584 2920
rect 7694 2812 7742 2920
rect 7852 2812 7900 2920
rect 8010 2812 8058 2920
rect 8168 2812 8216 2920
rect 8326 2812 8374 2920
rect 8484 2812 8532 2920
rect 8642 2812 8690 2920
rect 8800 2812 8848 2920
rect 8958 2812 9006 2920
rect 9116 2812 9164 2920
rect 9274 2812 9322 2920
rect 9432 2812 9480 2920
rect 9590 2812 9638 2920
rect 9748 2812 9796 2920
rect 9906 2812 9954 2920
rect 10064 2812 10112 2920
rect 10222 2812 10270 2920
rect 10380 2812 10428 2920
rect 10538 2812 10586 2920
rect 10696 2812 10744 2920
rect 10854 2812 10902 2920
rect 11012 2812 11060 2920
rect 11170 2812 11218 2920
rect 11328 2812 11376 2920
rect 11486 2812 11534 2920
rect 11644 2812 11692 2920
rect 11802 2812 11850 2920
rect 11960 2812 12008 2920
rect 12118 2812 12166 2920
rect 12276 2812 12324 2920
rect 12434 2812 12482 2920
rect 12592 2812 12640 2920
rect 12744 2812 12798 2920
rect 98 2804 172 2812
rect 98 2802 110 2804
rect 162 2802 172 2804
rect 98 2024 108 2802
rect 164 2024 172 2802
rect 98 2022 110 2024
rect 162 2022 172 2024
rect 98 2014 172 2022
rect 256 2802 328 2812
rect 256 2020 266 2802
rect 322 2020 328 2802
rect 110 1902 158 2014
rect 256 2010 328 2020
rect 412 2804 488 2812
rect 412 2802 426 2804
rect 412 2020 422 2802
rect 478 2020 488 2804
rect 412 2010 488 2020
rect 572 2802 644 2812
rect 572 2020 582 2802
rect 638 2020 644 2802
rect 572 2010 644 2020
rect 728 2804 804 2812
rect 728 2802 742 2804
rect 728 2020 738 2802
rect 794 2020 804 2804
rect 728 2010 804 2020
rect 888 2802 960 2812
rect 888 2020 898 2802
rect 954 2020 960 2802
rect 888 2010 960 2020
rect 1044 2804 1120 2812
rect 1044 2802 1058 2804
rect 1044 2020 1054 2802
rect 1110 2020 1120 2804
rect 1044 2010 1120 2020
rect 1204 2802 1276 2812
rect 1204 2020 1214 2802
rect 1270 2020 1276 2802
rect 1204 2010 1276 2020
rect 1360 2804 1436 2812
rect 1360 2802 1374 2804
rect 1360 2020 1370 2802
rect 1426 2020 1436 2804
rect 1360 2010 1436 2020
rect 1520 2802 1592 2812
rect 1520 2020 1530 2802
rect 1586 2020 1592 2802
rect 1520 2010 1592 2020
rect 1676 2804 1752 2812
rect 1676 2802 1690 2804
rect 1676 2020 1686 2802
rect 1742 2020 1752 2804
rect 1676 2010 1752 2020
rect 1836 2802 1908 2812
rect 1836 2020 1846 2802
rect 1902 2020 1908 2802
rect 1836 2010 1908 2020
rect 1992 2804 2068 2812
rect 1992 2802 2006 2804
rect 1992 2020 2002 2802
rect 2058 2020 2068 2804
rect 1992 2010 2068 2020
rect 2152 2802 2224 2812
rect 2152 2020 2162 2802
rect 2218 2020 2224 2802
rect 2152 2010 2224 2020
rect 2308 2804 2384 2812
rect 2308 2802 2322 2804
rect 2308 2020 2318 2802
rect 2374 2020 2384 2804
rect 2308 2010 2384 2020
rect 2468 2802 2540 2812
rect 2468 2020 2478 2802
rect 2534 2020 2540 2802
rect 2468 2010 2540 2020
rect 2624 2804 2700 2812
rect 2624 2802 2638 2804
rect 2624 2020 2634 2802
rect 2690 2020 2700 2804
rect 2624 2010 2700 2020
rect 2784 2802 2856 2812
rect 2784 2020 2794 2802
rect 2850 2020 2856 2802
rect 2784 2010 2856 2020
rect 2940 2804 3016 2812
rect 2940 2802 2954 2804
rect 2940 2020 2950 2802
rect 3006 2020 3016 2804
rect 2940 2010 3016 2020
rect 3100 2802 3172 2812
rect 3100 2020 3110 2802
rect 3166 2020 3172 2802
rect 3100 2010 3172 2020
rect 3256 2804 3332 2812
rect 3256 2802 3270 2804
rect 3256 2020 3266 2802
rect 3322 2020 3332 2804
rect 3256 2010 3332 2020
rect 3416 2802 3488 2812
rect 3416 2020 3426 2802
rect 3482 2020 3488 2802
rect 3416 2010 3488 2020
rect 3572 2804 3648 2812
rect 3572 2802 3586 2804
rect 3572 2020 3582 2802
rect 3638 2020 3648 2804
rect 3572 2010 3648 2020
rect 3732 2802 3804 2812
rect 3732 2020 3742 2802
rect 3798 2020 3804 2802
rect 3732 2010 3804 2020
rect 3888 2804 3964 2812
rect 3888 2802 3902 2804
rect 3888 2020 3898 2802
rect 3954 2020 3964 2804
rect 3888 2010 3964 2020
rect 4048 2802 4120 2812
rect 4048 2020 4058 2802
rect 4114 2020 4120 2802
rect 4048 2010 4120 2020
rect 4204 2804 4280 2812
rect 4204 2802 4218 2804
rect 4204 2020 4214 2802
rect 4270 2020 4280 2804
rect 4204 2010 4280 2020
rect 4364 2802 4436 2812
rect 4364 2020 4374 2802
rect 4430 2020 4436 2802
rect 4364 2010 4436 2020
rect 4520 2804 4596 2812
rect 4520 2802 4534 2804
rect 4520 2020 4530 2802
rect 4586 2020 4596 2804
rect 4520 2010 4596 2020
rect 4680 2802 4752 2812
rect 4680 2020 4690 2802
rect 4746 2020 4752 2802
rect 4680 2010 4752 2020
rect 4836 2804 4912 2812
rect 4836 2802 4850 2804
rect 4836 2020 4846 2802
rect 4902 2020 4912 2804
rect 4836 2010 4912 2020
rect 4996 2802 5068 2812
rect 4996 2020 5006 2802
rect 5062 2020 5068 2802
rect 4996 2010 5068 2020
rect 5152 2804 5228 2812
rect 5152 2802 5166 2804
rect 5152 2020 5162 2802
rect 5218 2020 5228 2804
rect 5152 2010 5228 2020
rect 5312 2802 5384 2812
rect 5312 2020 5322 2802
rect 5378 2020 5384 2802
rect 5312 2010 5384 2020
rect 5468 2804 5544 2812
rect 5468 2802 5482 2804
rect 5468 2020 5478 2802
rect 5534 2020 5544 2804
rect 5468 2010 5544 2020
rect 5628 2802 5700 2812
rect 5628 2020 5638 2802
rect 5694 2020 5700 2802
rect 5628 2010 5700 2020
rect 5784 2804 5860 2812
rect 5784 2802 5798 2804
rect 5784 2020 5794 2802
rect 5850 2020 5860 2804
rect 5784 2010 5860 2020
rect 5944 2802 6016 2812
rect 5944 2020 5954 2802
rect 6010 2020 6016 2802
rect 5944 2010 6016 2020
rect 6100 2804 6176 2812
rect 6100 2802 6114 2804
rect 6100 2020 6110 2802
rect 6166 2020 6176 2804
rect 6100 2010 6176 2020
rect 6260 2802 6332 2812
rect 6260 2020 6270 2802
rect 6326 2020 6332 2802
rect 6260 2010 6332 2020
rect 6416 2804 6492 2812
rect 6416 2802 6430 2804
rect 6416 2020 6426 2802
rect 6482 2020 6492 2804
rect 6416 2010 6492 2020
rect 6576 2802 6648 2812
rect 6576 2020 6586 2802
rect 6642 2020 6648 2802
rect 6576 2010 6648 2020
rect 6732 2804 6808 2812
rect 6732 2802 6746 2804
rect 6732 2020 6742 2802
rect 6798 2020 6808 2804
rect 6732 2010 6808 2020
rect 6892 2802 6964 2812
rect 6892 2020 6902 2802
rect 6958 2020 6964 2802
rect 6892 2010 6964 2020
rect 7048 2804 7124 2812
rect 7048 2802 7062 2804
rect 7048 2020 7058 2802
rect 7114 2020 7124 2804
rect 7048 2010 7124 2020
rect 7208 2802 7280 2812
rect 7208 2020 7218 2802
rect 7274 2020 7280 2802
rect 7208 2010 7280 2020
rect 7364 2804 7440 2812
rect 7364 2802 7378 2804
rect 7364 2020 7374 2802
rect 7430 2020 7440 2804
rect 7364 2010 7440 2020
rect 7524 2802 7596 2812
rect 7524 2020 7534 2802
rect 7590 2020 7596 2802
rect 7524 2010 7596 2020
rect 7680 2804 7756 2812
rect 7680 2802 7694 2804
rect 7680 2020 7690 2802
rect 7746 2020 7756 2804
rect 7680 2010 7756 2020
rect 7840 2802 7912 2812
rect 7840 2020 7850 2802
rect 7906 2020 7912 2802
rect 7840 2010 7912 2020
rect 7996 2804 8072 2812
rect 7996 2802 8010 2804
rect 7996 2020 8006 2802
rect 8062 2020 8072 2804
rect 7996 2010 8072 2020
rect 8156 2802 8228 2812
rect 8156 2020 8166 2802
rect 8222 2020 8228 2802
rect 8156 2010 8228 2020
rect 8312 2804 8388 2812
rect 8312 2802 8326 2804
rect 8312 2020 8322 2802
rect 8378 2020 8388 2804
rect 8312 2010 8388 2020
rect 8472 2802 8544 2812
rect 8472 2020 8482 2802
rect 8538 2020 8544 2802
rect 8472 2010 8544 2020
rect 8628 2804 8704 2812
rect 8628 2802 8642 2804
rect 8628 2020 8638 2802
rect 8694 2020 8704 2804
rect 8628 2010 8704 2020
rect 8788 2802 8860 2812
rect 8788 2020 8798 2802
rect 8854 2020 8860 2802
rect 8788 2010 8860 2020
rect 8944 2804 9020 2812
rect 8944 2802 8958 2804
rect 8944 2020 8954 2802
rect 9010 2020 9020 2804
rect 8944 2010 9020 2020
rect 9104 2802 9176 2812
rect 9104 2020 9114 2802
rect 9170 2020 9176 2802
rect 9104 2010 9176 2020
rect 9260 2804 9336 2812
rect 9260 2802 9274 2804
rect 9260 2020 9270 2802
rect 9326 2020 9336 2804
rect 9260 2010 9336 2020
rect 9420 2802 9492 2812
rect 9420 2020 9430 2802
rect 9486 2020 9492 2802
rect 9420 2010 9492 2020
rect 9576 2804 9652 2812
rect 9576 2802 9590 2804
rect 9576 2020 9586 2802
rect 9642 2020 9652 2804
rect 9576 2010 9652 2020
rect 9736 2802 9808 2812
rect 9736 2020 9746 2802
rect 9802 2020 9808 2802
rect 9736 2010 9808 2020
rect 9892 2804 9968 2812
rect 9892 2802 9906 2804
rect 9892 2020 9902 2802
rect 9958 2020 9968 2804
rect 9892 2010 9968 2020
rect 10052 2802 10124 2812
rect 10052 2020 10062 2802
rect 10118 2020 10124 2802
rect 10052 2010 10124 2020
rect 10208 2804 10284 2812
rect 10208 2802 10222 2804
rect 10208 2020 10218 2802
rect 10274 2020 10284 2804
rect 10208 2010 10284 2020
rect 10368 2802 10440 2812
rect 10368 2020 10378 2802
rect 10434 2020 10440 2802
rect 10368 2010 10440 2020
rect 10524 2804 10600 2812
rect 10524 2802 10538 2804
rect 10524 2020 10534 2802
rect 10590 2020 10600 2804
rect 10524 2010 10600 2020
rect 10684 2802 10756 2812
rect 10684 2020 10694 2802
rect 10750 2020 10756 2802
rect 10684 2010 10756 2020
rect 10840 2804 10916 2812
rect 10840 2802 10854 2804
rect 10840 2020 10850 2802
rect 10906 2020 10916 2804
rect 10840 2010 10916 2020
rect 11000 2802 11072 2812
rect 11000 2020 11010 2802
rect 11066 2020 11072 2802
rect 11000 2010 11072 2020
rect 11156 2804 11232 2812
rect 11156 2802 11170 2804
rect 11156 2020 11166 2802
rect 11222 2020 11232 2804
rect 11156 2010 11232 2020
rect 11316 2802 11388 2812
rect 11316 2020 11326 2802
rect 11382 2020 11388 2802
rect 11316 2010 11388 2020
rect 11472 2804 11548 2812
rect 11472 2802 11486 2804
rect 11472 2020 11482 2802
rect 11538 2020 11548 2804
rect 11472 2010 11548 2020
rect 11632 2802 11704 2812
rect 11632 2020 11642 2802
rect 11698 2020 11704 2802
rect 11632 2010 11704 2020
rect 11788 2804 11864 2812
rect 11788 2802 11802 2804
rect 11788 2020 11798 2802
rect 11854 2020 11864 2804
rect 11788 2010 11864 2020
rect 11948 2802 12020 2812
rect 11948 2020 11958 2802
rect 12014 2020 12020 2802
rect 11948 2010 12020 2020
rect 12104 2804 12180 2812
rect 12104 2802 12118 2804
rect 12104 2020 12114 2802
rect 12170 2020 12180 2804
rect 12104 2010 12180 2020
rect 12264 2802 12336 2812
rect 12264 2020 12274 2802
rect 12330 2020 12336 2802
rect 12264 2010 12336 2020
rect 12420 2804 12496 2812
rect 12420 2802 12434 2804
rect 12420 2020 12430 2802
rect 12486 2020 12496 2804
rect 12420 2010 12496 2020
rect 12580 2802 12652 2812
rect 12580 2020 12590 2802
rect 12646 2020 12652 2802
rect 12580 2010 12652 2020
rect 12736 2804 12812 2812
rect 12736 2022 12744 2804
rect 12796 2802 12812 2804
rect 12736 2020 12746 2022
rect 12802 2020 12812 2802
rect 12736 2010 12812 2020
rect 268 1902 316 2010
rect 426 1902 474 2010
rect 584 1902 632 2010
rect 742 1902 790 2010
rect 900 1902 948 2010
rect 1058 1902 1106 2010
rect 1216 1902 1264 2010
rect 1374 1902 1422 2010
rect 1532 1902 1580 2010
rect 1690 1902 1738 2010
rect 1848 1902 1896 2010
rect 2006 1902 2054 2010
rect 2164 1902 2212 2010
rect 2322 1902 2370 2010
rect 2480 1902 2528 2010
rect 2638 1902 2686 2010
rect 2796 1902 2844 2010
rect 2954 1902 3002 2010
rect 3112 1902 3160 2010
rect 3270 1902 3318 2010
rect 3428 1902 3476 2010
rect 3586 1902 3634 2010
rect 3744 1902 3792 2010
rect 3902 1902 3950 2010
rect 4060 1902 4108 2010
rect 4218 1902 4266 2010
rect 4376 1902 4424 2010
rect 4534 1902 4582 2010
rect 4692 1902 4740 2010
rect 4850 1902 4898 2010
rect 5008 1902 5056 2010
rect 5166 1902 5214 2010
rect 5324 1902 5372 2010
rect 5482 1902 5530 2010
rect 5640 1902 5688 2010
rect 5798 1902 5846 2010
rect 5956 1902 6004 2010
rect 6114 1902 6162 2010
rect 6272 1902 6320 2010
rect 6430 1902 6478 2010
rect 6588 1902 6636 2010
rect 6746 1902 6794 2010
rect 6904 1902 6952 2010
rect 7062 1902 7110 2010
rect 7220 1902 7268 2010
rect 7378 1902 7426 2010
rect 7536 1902 7584 2010
rect 7694 1902 7742 2010
rect 7852 1902 7900 2010
rect 8010 1902 8058 2010
rect 8168 1902 8216 2010
rect 8326 1902 8374 2010
rect 8484 1902 8532 2010
rect 8642 1902 8690 2010
rect 8800 1902 8848 2010
rect 8958 1902 9006 2010
rect 9116 1902 9164 2010
rect 9274 1902 9322 2010
rect 9432 1902 9480 2010
rect 9590 1902 9638 2010
rect 9748 1902 9796 2010
rect 9906 1902 9954 2010
rect 10064 1902 10112 2010
rect 10222 1902 10270 2010
rect 10380 1902 10428 2010
rect 10538 1902 10586 2010
rect 10696 1902 10744 2010
rect 10854 1902 10902 2010
rect 11012 1902 11060 2010
rect 11170 1902 11218 2010
rect 11328 1902 11376 2010
rect 11486 1902 11534 2010
rect 11644 1902 11692 2010
rect 11802 1902 11850 2010
rect 11960 1902 12008 2010
rect 12118 1902 12166 2010
rect 12276 1902 12324 2010
rect 12434 1902 12482 2010
rect 12592 1902 12640 2010
rect 12744 1902 12798 2010
rect 98 1894 172 1902
rect 98 1892 110 1894
rect 162 1892 172 1894
rect 98 1114 108 1892
rect 164 1114 172 1892
rect 98 1112 110 1114
rect 162 1112 172 1114
rect 98 1104 172 1112
rect 256 1892 328 1902
rect 256 1110 266 1892
rect 322 1110 328 1892
rect 110 992 158 1104
rect 256 1100 328 1110
rect 412 1894 488 1902
rect 412 1892 426 1894
rect 412 1110 422 1892
rect 478 1110 488 1894
rect 412 1100 488 1110
rect 572 1892 644 1902
rect 572 1110 582 1892
rect 638 1110 644 1892
rect 572 1100 644 1110
rect 728 1894 804 1902
rect 728 1892 742 1894
rect 728 1110 738 1892
rect 794 1110 804 1894
rect 728 1100 804 1110
rect 888 1892 960 1902
rect 888 1110 898 1892
rect 954 1110 960 1892
rect 888 1100 960 1110
rect 1044 1894 1120 1902
rect 1044 1892 1058 1894
rect 1044 1110 1054 1892
rect 1110 1110 1120 1894
rect 1044 1100 1120 1110
rect 1204 1892 1276 1902
rect 1204 1110 1214 1892
rect 1270 1110 1276 1892
rect 1204 1100 1276 1110
rect 1360 1894 1436 1902
rect 1360 1892 1374 1894
rect 1360 1110 1370 1892
rect 1426 1110 1436 1894
rect 1360 1100 1436 1110
rect 1520 1892 1592 1902
rect 1520 1110 1530 1892
rect 1586 1110 1592 1892
rect 1520 1100 1592 1110
rect 1676 1894 1752 1902
rect 1676 1892 1690 1894
rect 1676 1110 1686 1892
rect 1742 1110 1752 1894
rect 1676 1100 1752 1110
rect 1836 1892 1908 1902
rect 1836 1110 1846 1892
rect 1902 1110 1908 1892
rect 1836 1100 1908 1110
rect 1992 1894 2068 1902
rect 1992 1892 2006 1894
rect 1992 1110 2002 1892
rect 2058 1110 2068 1894
rect 1992 1100 2068 1110
rect 2152 1892 2224 1902
rect 2152 1110 2162 1892
rect 2218 1110 2224 1892
rect 2152 1100 2224 1110
rect 2308 1894 2384 1902
rect 2308 1892 2322 1894
rect 2308 1110 2318 1892
rect 2374 1110 2384 1894
rect 2308 1100 2384 1110
rect 2468 1892 2540 1902
rect 2468 1110 2478 1892
rect 2534 1110 2540 1892
rect 2468 1100 2540 1110
rect 2624 1894 2700 1902
rect 2624 1892 2638 1894
rect 2624 1110 2634 1892
rect 2690 1110 2700 1894
rect 2624 1100 2700 1110
rect 2784 1892 2856 1902
rect 2784 1110 2794 1892
rect 2850 1110 2856 1892
rect 2784 1100 2856 1110
rect 2940 1894 3016 1902
rect 2940 1892 2954 1894
rect 2940 1110 2950 1892
rect 3006 1110 3016 1894
rect 2940 1100 3016 1110
rect 3100 1892 3172 1902
rect 3100 1110 3110 1892
rect 3166 1110 3172 1892
rect 3100 1100 3172 1110
rect 3256 1894 3332 1902
rect 3256 1892 3270 1894
rect 3256 1110 3266 1892
rect 3322 1110 3332 1894
rect 3256 1100 3332 1110
rect 3416 1892 3488 1902
rect 3416 1110 3426 1892
rect 3482 1110 3488 1892
rect 3416 1100 3488 1110
rect 3572 1894 3648 1902
rect 3572 1892 3586 1894
rect 3572 1110 3582 1892
rect 3638 1110 3648 1894
rect 3572 1100 3648 1110
rect 3732 1892 3804 1902
rect 3732 1110 3742 1892
rect 3798 1110 3804 1892
rect 3732 1100 3804 1110
rect 3888 1894 3964 1902
rect 3888 1892 3902 1894
rect 3888 1110 3898 1892
rect 3954 1110 3964 1894
rect 3888 1100 3964 1110
rect 4048 1892 4120 1902
rect 4048 1110 4058 1892
rect 4114 1110 4120 1892
rect 4048 1100 4120 1110
rect 4204 1894 4280 1902
rect 4204 1892 4218 1894
rect 4204 1110 4214 1892
rect 4270 1110 4280 1894
rect 4204 1100 4280 1110
rect 4364 1892 4436 1902
rect 4364 1110 4374 1892
rect 4430 1110 4436 1892
rect 4364 1100 4436 1110
rect 4520 1894 4596 1902
rect 4520 1892 4534 1894
rect 4520 1110 4530 1892
rect 4586 1110 4596 1894
rect 4520 1100 4596 1110
rect 4680 1892 4752 1902
rect 4680 1110 4690 1892
rect 4746 1110 4752 1892
rect 4680 1100 4752 1110
rect 4836 1894 4912 1902
rect 4836 1892 4850 1894
rect 4836 1110 4846 1892
rect 4902 1110 4912 1894
rect 4836 1100 4912 1110
rect 4996 1892 5068 1902
rect 4996 1110 5006 1892
rect 5062 1110 5068 1892
rect 4996 1100 5068 1110
rect 5152 1894 5228 1902
rect 5152 1892 5166 1894
rect 5152 1110 5162 1892
rect 5218 1110 5228 1894
rect 5152 1100 5228 1110
rect 5312 1892 5384 1902
rect 5312 1110 5322 1892
rect 5378 1110 5384 1892
rect 5312 1100 5384 1110
rect 5468 1894 5544 1902
rect 5468 1892 5482 1894
rect 5468 1110 5478 1892
rect 5534 1110 5544 1894
rect 5468 1100 5544 1110
rect 5628 1892 5700 1902
rect 5628 1110 5638 1892
rect 5694 1110 5700 1892
rect 5628 1100 5700 1110
rect 5784 1894 5860 1902
rect 5784 1892 5798 1894
rect 5784 1110 5794 1892
rect 5850 1110 5860 1894
rect 5784 1100 5860 1110
rect 5944 1892 6016 1902
rect 5944 1110 5954 1892
rect 6010 1110 6016 1892
rect 5944 1100 6016 1110
rect 6100 1894 6176 1902
rect 6100 1892 6114 1894
rect 6100 1110 6110 1892
rect 6166 1110 6176 1894
rect 6100 1100 6176 1110
rect 6260 1892 6332 1902
rect 6260 1110 6270 1892
rect 6326 1110 6332 1892
rect 6260 1100 6332 1110
rect 6416 1894 6492 1902
rect 6416 1892 6430 1894
rect 6416 1110 6426 1892
rect 6482 1110 6492 1894
rect 6416 1100 6492 1110
rect 6576 1892 6648 1902
rect 6576 1110 6586 1892
rect 6642 1110 6648 1892
rect 6576 1100 6648 1110
rect 6732 1894 6808 1902
rect 6732 1892 6746 1894
rect 6732 1110 6742 1892
rect 6798 1110 6808 1894
rect 6732 1100 6808 1110
rect 6892 1892 6964 1902
rect 6892 1110 6902 1892
rect 6958 1110 6964 1892
rect 6892 1100 6964 1110
rect 7048 1894 7124 1902
rect 7048 1892 7062 1894
rect 7048 1110 7058 1892
rect 7114 1110 7124 1894
rect 7048 1100 7124 1110
rect 7208 1892 7280 1902
rect 7208 1110 7218 1892
rect 7274 1110 7280 1892
rect 7208 1100 7280 1110
rect 7364 1894 7440 1902
rect 7364 1892 7378 1894
rect 7364 1110 7374 1892
rect 7430 1110 7440 1894
rect 7364 1100 7440 1110
rect 7524 1892 7596 1902
rect 7524 1110 7534 1892
rect 7590 1110 7596 1892
rect 7524 1100 7596 1110
rect 7680 1894 7756 1902
rect 7680 1892 7694 1894
rect 7680 1110 7690 1892
rect 7746 1110 7756 1894
rect 7680 1100 7756 1110
rect 7840 1892 7912 1902
rect 7840 1110 7850 1892
rect 7906 1110 7912 1892
rect 7840 1100 7912 1110
rect 7996 1894 8072 1902
rect 7996 1892 8010 1894
rect 7996 1110 8006 1892
rect 8062 1110 8072 1894
rect 7996 1100 8072 1110
rect 8156 1892 8228 1902
rect 8156 1110 8166 1892
rect 8222 1110 8228 1892
rect 8156 1100 8228 1110
rect 8312 1894 8388 1902
rect 8312 1892 8326 1894
rect 8312 1110 8322 1892
rect 8378 1110 8388 1894
rect 8312 1100 8388 1110
rect 8472 1892 8544 1902
rect 8472 1110 8482 1892
rect 8538 1110 8544 1892
rect 8472 1100 8544 1110
rect 8628 1894 8704 1902
rect 8628 1892 8642 1894
rect 8628 1110 8638 1892
rect 8694 1110 8704 1894
rect 8628 1100 8704 1110
rect 8788 1892 8860 1902
rect 8788 1110 8798 1892
rect 8854 1110 8860 1892
rect 8788 1100 8860 1110
rect 8944 1894 9020 1902
rect 8944 1892 8958 1894
rect 8944 1110 8954 1892
rect 9010 1110 9020 1894
rect 8944 1100 9020 1110
rect 9104 1892 9176 1902
rect 9104 1110 9114 1892
rect 9170 1110 9176 1892
rect 9104 1100 9176 1110
rect 9260 1894 9336 1902
rect 9260 1892 9274 1894
rect 9260 1110 9270 1892
rect 9326 1110 9336 1894
rect 9260 1100 9336 1110
rect 9420 1892 9492 1902
rect 9420 1110 9430 1892
rect 9486 1110 9492 1892
rect 9420 1100 9492 1110
rect 9576 1894 9652 1902
rect 9576 1892 9590 1894
rect 9576 1110 9586 1892
rect 9642 1110 9652 1894
rect 9576 1100 9652 1110
rect 9736 1892 9808 1902
rect 9736 1110 9746 1892
rect 9802 1110 9808 1892
rect 9736 1100 9808 1110
rect 9892 1894 9968 1902
rect 9892 1892 9906 1894
rect 9892 1110 9902 1892
rect 9958 1110 9968 1894
rect 9892 1100 9968 1110
rect 10052 1892 10124 1902
rect 10052 1110 10062 1892
rect 10118 1110 10124 1892
rect 10052 1100 10124 1110
rect 10208 1894 10284 1902
rect 10208 1892 10222 1894
rect 10208 1110 10218 1892
rect 10274 1110 10284 1894
rect 10208 1100 10284 1110
rect 10368 1892 10440 1902
rect 10368 1110 10378 1892
rect 10434 1110 10440 1892
rect 10368 1100 10440 1110
rect 10524 1894 10600 1902
rect 10524 1892 10538 1894
rect 10524 1110 10534 1892
rect 10590 1110 10600 1894
rect 10524 1100 10600 1110
rect 10684 1892 10756 1902
rect 10684 1110 10694 1892
rect 10750 1110 10756 1892
rect 10684 1100 10756 1110
rect 10840 1894 10916 1902
rect 10840 1892 10854 1894
rect 10840 1110 10850 1892
rect 10906 1110 10916 1894
rect 10840 1100 10916 1110
rect 11000 1892 11072 1902
rect 11000 1110 11010 1892
rect 11066 1110 11072 1892
rect 11000 1100 11072 1110
rect 11156 1894 11232 1902
rect 11156 1892 11170 1894
rect 11156 1110 11166 1892
rect 11222 1110 11232 1894
rect 11156 1100 11232 1110
rect 11316 1892 11388 1902
rect 11316 1110 11326 1892
rect 11382 1110 11388 1892
rect 11316 1100 11388 1110
rect 11472 1894 11548 1902
rect 11472 1892 11486 1894
rect 11472 1110 11482 1892
rect 11538 1110 11548 1894
rect 11472 1100 11548 1110
rect 11632 1892 11704 1902
rect 11632 1110 11642 1892
rect 11698 1110 11704 1892
rect 11632 1100 11704 1110
rect 11788 1894 11864 1902
rect 11788 1892 11802 1894
rect 11788 1110 11798 1892
rect 11854 1110 11864 1894
rect 11788 1100 11864 1110
rect 11948 1892 12020 1902
rect 11948 1110 11958 1892
rect 12014 1110 12020 1892
rect 11948 1100 12020 1110
rect 12104 1894 12180 1902
rect 12104 1892 12118 1894
rect 12104 1110 12114 1892
rect 12170 1110 12180 1894
rect 12104 1100 12180 1110
rect 12264 1892 12336 1902
rect 12264 1110 12274 1892
rect 12330 1110 12336 1892
rect 12264 1100 12336 1110
rect 12420 1894 12496 1902
rect 12420 1892 12434 1894
rect 12420 1110 12430 1892
rect 12486 1110 12496 1894
rect 12420 1100 12496 1110
rect 12580 1892 12652 1902
rect 12580 1110 12590 1892
rect 12646 1110 12652 1892
rect 12580 1100 12652 1110
rect 12736 1894 12812 1902
rect 12736 1112 12744 1894
rect 12796 1892 12812 1894
rect 12736 1110 12746 1112
rect 12802 1110 12812 1892
rect 12736 1100 12812 1110
rect 268 992 316 1100
rect 426 992 474 1100
rect 584 992 632 1100
rect 742 992 790 1100
rect 900 992 948 1100
rect 1058 992 1106 1100
rect 1216 992 1264 1100
rect 1374 992 1422 1100
rect 1532 992 1580 1100
rect 1690 992 1738 1100
rect 1848 992 1896 1100
rect 2006 992 2054 1100
rect 2164 992 2212 1100
rect 2322 992 2370 1100
rect 2480 992 2528 1100
rect 2638 992 2686 1100
rect 2796 992 2844 1100
rect 2954 992 3002 1100
rect 3112 992 3160 1100
rect 3270 992 3318 1100
rect 3428 992 3476 1100
rect 3586 992 3634 1100
rect 3744 992 3792 1100
rect 3902 992 3950 1100
rect 4060 992 4108 1100
rect 4218 992 4266 1100
rect 4376 992 4424 1100
rect 4534 992 4582 1100
rect 4692 992 4740 1100
rect 4850 992 4898 1100
rect 5008 992 5056 1100
rect 5166 992 5214 1100
rect 5324 992 5372 1100
rect 5482 992 5530 1100
rect 5640 992 5688 1100
rect 5798 992 5846 1100
rect 5956 992 6004 1100
rect 6114 992 6162 1100
rect 6272 992 6320 1100
rect 6430 992 6478 1100
rect 6588 992 6636 1100
rect 6746 992 6794 1100
rect 6904 992 6952 1100
rect 7062 992 7110 1100
rect 7220 992 7268 1100
rect 7378 992 7426 1100
rect 7536 992 7584 1100
rect 7694 992 7742 1100
rect 7852 992 7900 1100
rect 8010 992 8058 1100
rect 8168 992 8216 1100
rect 8326 992 8374 1100
rect 8484 992 8532 1100
rect 8642 992 8690 1100
rect 8800 992 8848 1100
rect 8958 992 9006 1100
rect 9116 992 9164 1100
rect 9274 992 9322 1100
rect 9432 992 9480 1100
rect 9590 992 9638 1100
rect 9748 992 9796 1100
rect 9906 992 9954 1100
rect 10064 992 10112 1100
rect 10222 992 10270 1100
rect 10380 992 10428 1100
rect 10538 992 10586 1100
rect 10696 992 10744 1100
rect 10854 992 10902 1100
rect 11012 992 11060 1100
rect 11170 992 11218 1100
rect 11328 992 11376 1100
rect 11486 992 11534 1100
rect 11644 992 11692 1100
rect 11802 992 11850 1100
rect 11960 992 12008 1100
rect 12118 992 12166 1100
rect 12276 992 12324 1100
rect 12434 992 12482 1100
rect 12592 992 12640 1100
rect 12744 992 12798 1100
rect 98 984 172 992
rect 98 982 110 984
rect 162 982 172 984
rect 98 204 108 982
rect 164 204 172 982
rect 98 202 110 204
rect 162 202 172 204
rect 98 194 172 202
rect 256 982 328 992
rect 256 200 266 982
rect 322 200 328 982
rect 110 -66 158 194
rect 256 190 328 200
rect 412 984 488 992
rect 412 982 426 984
rect 412 200 422 982
rect 478 200 488 984
rect 412 190 488 200
rect 572 982 644 992
rect 572 200 582 982
rect 638 200 644 982
rect 572 190 644 200
rect 728 984 804 992
rect 728 982 742 984
rect 728 200 738 982
rect 794 200 804 984
rect 728 190 804 200
rect 888 982 960 992
rect 888 200 898 982
rect 954 200 960 982
rect 888 190 960 200
rect 1044 984 1120 992
rect 1044 982 1058 984
rect 1044 200 1054 982
rect 1110 200 1120 984
rect 1044 190 1120 200
rect 1204 982 1276 992
rect 1204 200 1214 982
rect 1270 200 1276 982
rect 1204 190 1276 200
rect 1360 984 1436 992
rect 1360 982 1374 984
rect 1360 200 1370 982
rect 1426 200 1436 984
rect 1360 190 1436 200
rect 1520 982 1592 992
rect 1520 200 1530 982
rect 1586 200 1592 982
rect 1520 190 1592 200
rect 1676 984 1752 992
rect 1676 982 1690 984
rect 1676 200 1686 982
rect 1742 200 1752 984
rect 1676 190 1752 200
rect 1836 982 1908 992
rect 1836 200 1846 982
rect 1902 200 1908 982
rect 1836 190 1908 200
rect 1992 984 2068 992
rect 1992 982 2006 984
rect 1992 200 2002 982
rect 2058 200 2068 984
rect 1992 190 2068 200
rect 2152 982 2224 992
rect 2152 200 2162 982
rect 2218 200 2224 982
rect 2152 190 2224 200
rect 2308 984 2384 992
rect 2308 982 2322 984
rect 2308 200 2318 982
rect 2374 200 2384 984
rect 2308 190 2384 200
rect 2468 982 2540 992
rect 2468 200 2478 982
rect 2534 200 2540 982
rect 2468 190 2540 200
rect 2624 984 2700 992
rect 2624 982 2638 984
rect 2624 200 2634 982
rect 2690 200 2700 984
rect 2624 190 2700 200
rect 2784 982 2856 992
rect 2784 200 2794 982
rect 2850 200 2856 982
rect 2784 190 2856 200
rect 2940 984 3016 992
rect 2940 982 2954 984
rect 2940 200 2950 982
rect 3006 200 3016 984
rect 2940 190 3016 200
rect 3100 982 3172 992
rect 3100 200 3110 982
rect 3166 200 3172 982
rect 3100 190 3172 200
rect 3256 984 3332 992
rect 3256 982 3270 984
rect 3256 200 3266 982
rect 3322 200 3332 984
rect 3256 190 3332 200
rect 3416 982 3488 992
rect 3416 200 3426 982
rect 3482 200 3488 982
rect 3416 190 3488 200
rect 3572 984 3648 992
rect 3572 982 3586 984
rect 3572 200 3582 982
rect 3638 200 3648 984
rect 3572 190 3648 200
rect 3732 982 3804 992
rect 3732 200 3742 982
rect 3798 200 3804 982
rect 3732 190 3804 200
rect 3888 984 3964 992
rect 3888 982 3902 984
rect 3888 200 3898 982
rect 3954 200 3964 984
rect 3888 190 3964 200
rect 4048 982 4120 992
rect 4048 200 4058 982
rect 4114 200 4120 982
rect 4048 190 4120 200
rect 4204 984 4280 992
rect 4204 982 4218 984
rect 4204 200 4214 982
rect 4270 200 4280 984
rect 4204 190 4280 200
rect 4364 982 4436 992
rect 4364 200 4374 982
rect 4430 200 4436 982
rect 4364 190 4436 200
rect 4520 984 4596 992
rect 4520 982 4534 984
rect 4520 200 4530 982
rect 4586 200 4596 984
rect 4520 190 4596 200
rect 4680 982 4752 992
rect 4680 200 4690 982
rect 4746 200 4752 982
rect 4680 190 4752 200
rect 4836 984 4912 992
rect 4836 982 4850 984
rect 4836 200 4846 982
rect 4902 200 4912 984
rect 4836 190 4912 200
rect 4996 982 5068 992
rect 4996 200 5006 982
rect 5062 200 5068 982
rect 4996 190 5068 200
rect 5152 984 5228 992
rect 5152 982 5166 984
rect 5152 200 5162 982
rect 5218 200 5228 984
rect 5152 190 5228 200
rect 5312 982 5384 992
rect 5312 200 5322 982
rect 5378 200 5384 982
rect 5312 190 5384 200
rect 5468 984 5544 992
rect 5468 982 5482 984
rect 5468 200 5478 982
rect 5534 200 5544 984
rect 5468 190 5544 200
rect 5628 982 5700 992
rect 5628 200 5638 982
rect 5694 200 5700 982
rect 5628 190 5700 200
rect 5784 984 5860 992
rect 5784 982 5798 984
rect 5784 200 5794 982
rect 5850 200 5860 984
rect 5784 190 5860 200
rect 5944 982 6016 992
rect 5944 200 5954 982
rect 6010 200 6016 982
rect 5944 190 6016 200
rect 6100 984 6176 992
rect 6100 982 6114 984
rect 6100 200 6110 982
rect 6166 200 6176 984
rect 6100 190 6176 200
rect 6260 982 6332 992
rect 6260 200 6270 982
rect 6326 200 6332 982
rect 6260 190 6332 200
rect 6416 984 6492 992
rect 6416 982 6430 984
rect 6416 200 6426 982
rect 6482 200 6492 984
rect 6416 190 6492 200
rect 6576 982 6648 992
rect 6576 200 6586 982
rect 6642 200 6648 982
rect 6576 190 6648 200
rect 6732 984 6808 992
rect 6732 982 6746 984
rect 6732 200 6742 982
rect 6798 200 6808 984
rect 6732 190 6808 200
rect 6892 982 6964 992
rect 6892 200 6902 982
rect 6958 200 6964 982
rect 6892 190 6964 200
rect 7048 984 7124 992
rect 7048 982 7062 984
rect 7048 200 7058 982
rect 7114 200 7124 984
rect 7048 190 7124 200
rect 7208 982 7280 992
rect 7208 200 7218 982
rect 7274 200 7280 982
rect 7208 190 7280 200
rect 7364 984 7440 992
rect 7364 982 7378 984
rect 7364 200 7374 982
rect 7430 200 7440 984
rect 7364 190 7440 200
rect 7524 982 7596 992
rect 7524 200 7534 982
rect 7590 200 7596 982
rect 7524 190 7596 200
rect 7680 984 7756 992
rect 7680 982 7694 984
rect 7680 200 7690 982
rect 7746 200 7756 984
rect 7680 190 7756 200
rect 7840 982 7912 992
rect 7840 200 7850 982
rect 7906 200 7912 982
rect 7840 190 7912 200
rect 7996 984 8072 992
rect 7996 982 8010 984
rect 7996 200 8006 982
rect 8062 200 8072 984
rect 7996 190 8072 200
rect 8156 982 8228 992
rect 8156 200 8166 982
rect 8222 200 8228 982
rect 8156 190 8228 200
rect 8312 984 8388 992
rect 8312 982 8326 984
rect 8312 200 8322 982
rect 8378 200 8388 984
rect 8312 190 8388 200
rect 8472 982 8544 992
rect 8472 200 8482 982
rect 8538 200 8544 982
rect 8472 190 8544 200
rect 8628 984 8704 992
rect 8628 982 8642 984
rect 8628 200 8638 982
rect 8694 200 8704 984
rect 8628 190 8704 200
rect 8788 982 8860 992
rect 8788 200 8798 982
rect 8854 200 8860 982
rect 8788 190 8860 200
rect 8944 984 9020 992
rect 8944 982 8958 984
rect 8944 200 8954 982
rect 9010 200 9020 984
rect 8944 190 9020 200
rect 9104 982 9176 992
rect 9104 200 9114 982
rect 9170 200 9176 982
rect 9104 190 9176 200
rect 9260 984 9336 992
rect 9260 982 9274 984
rect 9260 200 9270 982
rect 9326 200 9336 984
rect 9260 190 9336 200
rect 9420 982 9492 992
rect 9420 200 9430 982
rect 9486 200 9492 982
rect 9420 190 9492 200
rect 9576 984 9652 992
rect 9576 982 9590 984
rect 9576 200 9586 982
rect 9642 200 9652 984
rect 9576 190 9652 200
rect 9736 982 9808 992
rect 9736 200 9746 982
rect 9802 200 9808 982
rect 9736 190 9808 200
rect 9892 984 9968 992
rect 9892 982 9906 984
rect 9892 200 9902 982
rect 9958 200 9968 984
rect 9892 190 9968 200
rect 10052 982 10124 992
rect 10052 200 10062 982
rect 10118 200 10124 982
rect 10052 190 10124 200
rect 10208 984 10284 992
rect 10208 982 10222 984
rect 10208 200 10218 982
rect 10274 200 10284 984
rect 10208 190 10284 200
rect 10368 982 10440 992
rect 10368 200 10378 982
rect 10434 200 10440 982
rect 10368 190 10440 200
rect 10524 984 10600 992
rect 10524 982 10538 984
rect 10524 200 10534 982
rect 10590 200 10600 984
rect 10524 190 10600 200
rect 10684 982 10756 992
rect 10684 200 10694 982
rect 10750 200 10756 982
rect 10684 190 10756 200
rect 10840 984 10916 992
rect 10840 982 10854 984
rect 10840 200 10850 982
rect 10906 200 10916 984
rect 10840 190 10916 200
rect 11000 982 11072 992
rect 11000 200 11010 982
rect 11066 200 11072 982
rect 11000 190 11072 200
rect 11156 984 11232 992
rect 11156 982 11170 984
rect 11156 200 11166 982
rect 11222 200 11232 984
rect 11156 190 11232 200
rect 11316 982 11388 992
rect 11316 200 11326 982
rect 11382 200 11388 982
rect 11316 190 11388 200
rect 11472 984 11548 992
rect 11472 982 11486 984
rect 11472 200 11482 982
rect 11538 200 11548 984
rect 11472 190 11548 200
rect 11632 982 11704 992
rect 11632 200 11642 982
rect 11698 200 11704 982
rect 11632 190 11704 200
rect 11788 984 11864 992
rect 11788 982 11802 984
rect 11788 200 11798 982
rect 11854 200 11864 984
rect 11788 190 11864 200
rect 11948 982 12020 992
rect 11948 200 11958 982
rect 12014 200 12020 982
rect 11948 190 12020 200
rect 12104 984 12180 992
rect 12104 982 12118 984
rect 12104 200 12114 982
rect 12170 200 12180 984
rect 12104 190 12180 200
rect 12264 982 12336 992
rect 12264 200 12274 982
rect 12330 200 12336 982
rect 12264 190 12336 200
rect 12420 984 12496 992
rect 12420 982 12434 984
rect 12420 200 12430 982
rect 12486 200 12496 984
rect 12420 190 12496 200
rect 12580 982 12652 992
rect 12580 200 12590 982
rect 12646 200 12652 982
rect 12580 190 12652 200
rect 12736 984 12812 992
rect 12736 202 12744 984
rect 12796 982 12812 984
rect 12736 200 12746 202
rect 12802 200 12812 982
rect 12736 190 12812 200
rect 268 32 316 190
rect 254 26 330 32
rect 254 -28 260 26
rect 324 -28 330 26
rect 254 -34 330 -28
rect 268 -66 316 -34
rect 426 -66 474 190
rect 584 32 632 190
rect 570 26 646 32
rect 570 -28 576 26
rect 640 -28 646 26
rect 570 -34 646 -28
rect 584 -66 632 -34
rect 742 -66 790 190
rect 900 32 948 190
rect 886 26 962 32
rect 886 -28 892 26
rect 956 -28 962 26
rect 886 -34 962 -28
rect 900 -66 948 -34
rect 1058 -66 1106 190
rect 1216 32 1264 190
rect 1202 26 1278 32
rect 1202 -28 1208 26
rect 1272 -28 1278 26
rect 1202 -34 1278 -28
rect 1216 -66 1264 -34
rect 1374 -66 1422 190
rect 1532 32 1580 190
rect 1518 26 1594 32
rect 1518 -28 1524 26
rect 1588 -28 1594 26
rect 1518 -34 1594 -28
rect 1532 -66 1580 -34
rect 1690 -66 1738 190
rect 1848 32 1896 190
rect 1834 26 1910 32
rect 1834 -28 1840 26
rect 1904 -28 1910 26
rect 1834 -34 1910 -28
rect 1848 -66 1896 -34
rect 2006 -66 2054 190
rect 2164 32 2212 190
rect 2150 26 2226 32
rect 2150 -28 2156 26
rect 2220 -28 2226 26
rect 2150 -34 2226 -28
rect 2164 -66 2212 -34
rect 2322 -66 2370 190
rect 2480 32 2528 190
rect 2466 26 2542 32
rect 2466 -28 2472 26
rect 2536 -28 2542 26
rect 2466 -34 2542 -28
rect 2480 -66 2528 -34
rect 2638 -66 2686 190
rect 2796 32 2844 190
rect 2782 26 2858 32
rect 2782 -28 2788 26
rect 2852 -28 2858 26
rect 2782 -34 2858 -28
rect 2796 -66 2844 -34
rect 2954 -66 3002 190
rect 3112 32 3160 190
rect 3098 26 3174 32
rect 3098 -28 3104 26
rect 3168 -28 3174 26
rect 3098 -34 3174 -28
rect 3112 -66 3160 -34
rect 3270 -66 3318 190
rect 3428 32 3476 190
rect 3414 26 3490 32
rect 3414 -28 3420 26
rect 3484 -28 3490 26
rect 3414 -34 3490 -28
rect 3428 -66 3476 -34
rect 3586 -66 3634 190
rect 3744 32 3792 190
rect 3730 26 3806 32
rect 3730 -28 3736 26
rect 3800 -28 3806 26
rect 3730 -34 3806 -28
rect 3744 -66 3792 -34
rect 3902 -66 3950 190
rect 4060 32 4108 190
rect 4046 26 4122 32
rect 4046 -28 4052 26
rect 4116 -28 4122 26
rect 4046 -34 4122 -28
rect 4060 -66 4108 -34
rect 4218 -66 4266 190
rect 4376 32 4424 190
rect 4362 26 4438 32
rect 4362 -28 4368 26
rect 4432 -28 4438 26
rect 4362 -34 4438 -28
rect 4376 -66 4424 -34
rect 4534 -66 4582 190
rect 4692 32 4740 190
rect 4678 26 4754 32
rect 4678 -28 4684 26
rect 4748 -28 4754 26
rect 4678 -34 4754 -28
rect 4692 -66 4740 -34
rect 4850 -66 4898 190
rect 5008 32 5056 190
rect 4994 26 5070 32
rect 4994 -28 5000 26
rect 5064 -28 5070 26
rect 4994 -34 5070 -28
rect 5008 -66 5056 -34
rect 5166 -66 5214 190
rect 5324 32 5372 190
rect 5310 26 5386 32
rect 5310 -28 5316 26
rect 5380 -28 5386 26
rect 5310 -34 5386 -28
rect 5324 -66 5372 -34
rect 5482 -66 5530 190
rect 5640 32 5688 190
rect 5626 26 5702 32
rect 5626 -28 5632 26
rect 5696 -28 5702 26
rect 5626 -34 5702 -28
rect 5640 -66 5688 -34
rect 5798 -66 5846 190
rect 5956 32 6004 190
rect 5942 26 6018 32
rect 5942 -28 5948 26
rect 6012 -28 6018 26
rect 5942 -34 6018 -28
rect 5956 -66 6004 -34
rect 6114 -66 6162 190
rect 6272 32 6320 190
rect 6258 26 6334 32
rect 6258 -28 6264 26
rect 6328 -28 6334 26
rect 6258 -34 6334 -28
rect 6272 -66 6320 -34
rect 6430 -66 6478 190
rect 6588 32 6636 190
rect 6574 26 6650 32
rect 6574 -28 6580 26
rect 6644 -28 6650 26
rect 6574 -34 6650 -28
rect 6588 -66 6636 -34
rect 6746 -66 6794 190
rect 6904 32 6952 190
rect 6890 26 6966 32
rect 6890 -28 6896 26
rect 6960 -28 6966 26
rect 6890 -34 6966 -28
rect 6904 -66 6952 -34
rect 7062 -66 7110 190
rect 7220 32 7268 190
rect 7206 26 7282 32
rect 7206 -28 7212 26
rect 7276 -28 7282 26
rect 7206 -34 7282 -28
rect 7220 -66 7268 -34
rect 7378 -66 7426 190
rect 7536 32 7584 190
rect 7522 26 7598 32
rect 7522 -28 7528 26
rect 7592 -28 7598 26
rect 7522 -34 7598 -28
rect 7536 -66 7584 -34
rect 7694 -66 7742 190
rect 7852 32 7900 190
rect 7838 26 7914 32
rect 7838 -28 7844 26
rect 7908 -28 7914 26
rect 7838 -34 7914 -28
rect 7852 -66 7900 -34
rect 8010 -66 8058 190
rect 8168 32 8216 190
rect 8154 26 8230 32
rect 8154 -28 8160 26
rect 8224 -28 8230 26
rect 8154 -34 8230 -28
rect 8168 -66 8216 -34
rect 8326 -66 8374 190
rect 8484 32 8532 190
rect 8470 26 8546 32
rect 8470 -28 8476 26
rect 8540 -28 8546 26
rect 8470 -34 8546 -28
rect 8484 -66 8532 -34
rect 8642 -66 8690 190
rect 8800 32 8848 190
rect 8786 26 8862 32
rect 8786 -28 8792 26
rect 8856 -28 8862 26
rect 8786 -34 8862 -28
rect 8800 -66 8848 -34
rect 8958 -66 9006 190
rect 9116 32 9164 190
rect 9102 26 9178 32
rect 9102 -28 9108 26
rect 9172 -28 9178 26
rect 9102 -34 9178 -28
rect 9116 -66 9164 -34
rect 9274 -66 9322 190
rect 9432 32 9480 190
rect 9418 26 9494 32
rect 9418 -28 9424 26
rect 9488 -28 9494 26
rect 9418 -34 9494 -28
rect 9432 -66 9480 -34
rect 9590 -66 9638 190
rect 9748 32 9796 190
rect 9734 26 9810 32
rect 9734 -28 9740 26
rect 9804 -28 9810 26
rect 9734 -34 9810 -28
rect 9748 -66 9796 -34
rect 9906 -66 9954 190
rect 10064 32 10112 190
rect 10050 26 10126 32
rect 10050 -28 10056 26
rect 10120 -28 10126 26
rect 10050 -34 10126 -28
rect 10064 -66 10112 -34
rect 10222 -66 10270 190
rect 10380 32 10428 190
rect 10366 26 10442 32
rect 10366 -28 10372 26
rect 10436 -28 10442 26
rect 10366 -34 10442 -28
rect 10380 -66 10428 -34
rect 10538 -66 10586 190
rect 10696 32 10744 190
rect 10682 26 10758 32
rect 10682 -28 10688 26
rect 10752 -28 10758 26
rect 10682 -34 10758 -28
rect 10696 -66 10744 -34
rect 10854 -66 10902 190
rect 11012 32 11060 190
rect 10998 26 11074 32
rect 10998 -28 11004 26
rect 11068 -28 11074 26
rect 10998 -34 11074 -28
rect 11012 -66 11060 -34
rect 11170 -66 11218 190
rect 11328 32 11376 190
rect 11314 26 11390 32
rect 11314 -28 11320 26
rect 11384 -28 11390 26
rect 11314 -34 11390 -28
rect 11328 -66 11376 -34
rect 11486 -66 11534 190
rect 11644 32 11692 190
rect 11630 26 11706 32
rect 11630 -28 11636 26
rect 11700 -28 11706 26
rect 11630 -34 11706 -28
rect 11644 -66 11692 -34
rect 11802 -66 11850 190
rect 11960 32 12008 190
rect 11946 26 12022 32
rect 11946 -28 11952 26
rect 12016 -28 12022 26
rect 11946 -34 12022 -28
rect 11960 -66 12008 -34
rect 12118 -66 12166 190
rect 12276 32 12324 190
rect 12262 26 12338 32
rect 12262 -28 12268 26
rect 12332 -28 12338 26
rect 12262 -34 12338 -28
rect 12276 -66 12324 -34
rect 12434 -66 12482 190
rect 12592 32 12640 190
rect 12578 26 12654 32
rect 12578 -28 12584 26
rect 12648 -28 12654 26
rect 12578 -34 12654 -28
rect 12592 -66 12640 -34
rect 12750 -66 12798 190
<< via2 >>
rect 108 3844 110 4622
rect 110 3844 162 4622
rect 162 3844 164 4622
rect 266 3840 268 4622
rect 268 3840 320 4622
rect 320 3840 322 4622
rect 422 3844 426 4622
rect 426 3844 478 4622
rect 422 3840 478 3844
rect 582 3840 584 4622
rect 584 3840 636 4622
rect 636 3840 638 4622
rect 738 3844 742 4622
rect 742 3844 794 4622
rect 738 3840 794 3844
rect 898 3840 900 4622
rect 900 3840 952 4622
rect 952 3840 954 4622
rect 1054 3844 1058 4622
rect 1058 3844 1110 4622
rect 1054 3840 1110 3844
rect 1214 3840 1216 4622
rect 1216 3840 1268 4622
rect 1268 3840 1270 4622
rect 1370 3844 1374 4622
rect 1374 3844 1426 4622
rect 1370 3840 1426 3844
rect 1530 3840 1532 4622
rect 1532 3840 1584 4622
rect 1584 3840 1586 4622
rect 1686 3844 1690 4622
rect 1690 3844 1742 4622
rect 1686 3840 1742 3844
rect 1846 3840 1848 4622
rect 1848 3840 1900 4622
rect 1900 3840 1902 4622
rect 2002 3844 2006 4622
rect 2006 3844 2058 4622
rect 2002 3840 2058 3844
rect 2162 3840 2164 4622
rect 2164 3840 2216 4622
rect 2216 3840 2218 4622
rect 2318 3844 2322 4622
rect 2322 3844 2374 4622
rect 2318 3840 2374 3844
rect 2478 3840 2480 4622
rect 2480 3840 2532 4622
rect 2532 3840 2534 4622
rect 2634 3844 2638 4622
rect 2638 3844 2690 4622
rect 2634 3840 2690 3844
rect 2794 3840 2796 4622
rect 2796 3840 2848 4622
rect 2848 3840 2850 4622
rect 2950 3844 2954 4622
rect 2954 3844 3006 4622
rect 2950 3840 3006 3844
rect 3110 3840 3112 4622
rect 3112 3840 3164 4622
rect 3164 3840 3166 4622
rect 3266 3844 3270 4622
rect 3270 3844 3322 4622
rect 3266 3840 3322 3844
rect 3426 3840 3428 4622
rect 3428 3840 3480 4622
rect 3480 3840 3482 4622
rect 3582 3844 3586 4622
rect 3586 3844 3638 4622
rect 3582 3840 3638 3844
rect 3742 3840 3744 4622
rect 3744 3840 3796 4622
rect 3796 3840 3798 4622
rect 3898 3844 3902 4622
rect 3902 3844 3954 4622
rect 3898 3840 3954 3844
rect 4058 3840 4060 4622
rect 4060 3840 4112 4622
rect 4112 3840 4114 4622
rect 4214 3844 4218 4622
rect 4218 3844 4270 4622
rect 4214 3840 4270 3844
rect 4374 3840 4376 4622
rect 4376 3840 4428 4622
rect 4428 3840 4430 4622
rect 4530 3844 4534 4622
rect 4534 3844 4586 4622
rect 4530 3840 4586 3844
rect 4690 3840 4692 4622
rect 4692 3840 4744 4622
rect 4744 3840 4746 4622
rect 4846 3844 4850 4622
rect 4850 3844 4902 4622
rect 4846 3840 4902 3844
rect 5006 3840 5008 4622
rect 5008 3840 5060 4622
rect 5060 3840 5062 4622
rect 5162 3844 5166 4622
rect 5166 3844 5218 4622
rect 5162 3840 5218 3844
rect 5322 3840 5324 4622
rect 5324 3840 5376 4622
rect 5376 3840 5378 4622
rect 5478 3844 5482 4622
rect 5482 3844 5534 4622
rect 5478 3840 5534 3844
rect 5638 3840 5640 4622
rect 5640 3840 5692 4622
rect 5692 3840 5694 4622
rect 5794 3844 5798 4622
rect 5798 3844 5850 4622
rect 5794 3840 5850 3844
rect 5954 3840 5956 4622
rect 5956 3840 6008 4622
rect 6008 3840 6010 4622
rect 6110 3844 6114 4622
rect 6114 3844 6166 4622
rect 6110 3840 6166 3844
rect 6270 3840 6272 4622
rect 6272 3840 6324 4622
rect 6324 3840 6326 4622
rect 6426 3844 6430 4622
rect 6430 3844 6482 4622
rect 6426 3840 6482 3844
rect 6586 3840 6588 4622
rect 6588 3840 6640 4622
rect 6640 3840 6642 4622
rect 6742 3844 6746 4622
rect 6746 3844 6798 4622
rect 6742 3840 6798 3844
rect 6902 3840 6904 4622
rect 6904 3840 6956 4622
rect 6956 3840 6958 4622
rect 7058 3844 7062 4622
rect 7062 3844 7114 4622
rect 7058 3840 7114 3844
rect 7218 3840 7220 4622
rect 7220 3840 7272 4622
rect 7272 3840 7274 4622
rect 7374 3844 7378 4622
rect 7378 3844 7430 4622
rect 7374 3840 7430 3844
rect 7534 3840 7536 4622
rect 7536 3840 7588 4622
rect 7588 3840 7590 4622
rect 7690 3844 7694 4622
rect 7694 3844 7746 4622
rect 7690 3840 7746 3844
rect 7850 3840 7852 4622
rect 7852 3840 7904 4622
rect 7904 3840 7906 4622
rect 8006 3844 8010 4622
rect 8010 3844 8062 4622
rect 8006 3840 8062 3844
rect 8166 3840 8168 4622
rect 8168 3840 8220 4622
rect 8220 3840 8222 4622
rect 8322 3844 8326 4622
rect 8326 3844 8378 4622
rect 8322 3840 8378 3844
rect 8482 3840 8484 4622
rect 8484 3840 8536 4622
rect 8536 3840 8538 4622
rect 8638 3844 8642 4622
rect 8642 3844 8694 4622
rect 8638 3840 8694 3844
rect 8798 3840 8800 4622
rect 8800 3840 8852 4622
rect 8852 3840 8854 4622
rect 8954 3844 8958 4622
rect 8958 3844 9010 4622
rect 8954 3840 9010 3844
rect 9114 3840 9116 4622
rect 9116 3840 9168 4622
rect 9168 3840 9170 4622
rect 9270 3844 9274 4622
rect 9274 3844 9326 4622
rect 9270 3840 9326 3844
rect 9430 3840 9432 4622
rect 9432 3840 9484 4622
rect 9484 3840 9486 4622
rect 9586 3844 9590 4622
rect 9590 3844 9642 4622
rect 9586 3840 9642 3844
rect 9746 3840 9748 4622
rect 9748 3840 9800 4622
rect 9800 3840 9802 4622
rect 9902 3844 9906 4622
rect 9906 3844 9958 4622
rect 9902 3840 9958 3844
rect 10062 3840 10064 4622
rect 10064 3840 10116 4622
rect 10116 3840 10118 4622
rect 10218 3844 10222 4622
rect 10222 3844 10274 4622
rect 10218 3840 10274 3844
rect 10378 3840 10380 4622
rect 10380 3840 10432 4622
rect 10432 3840 10434 4622
rect 10534 3844 10538 4622
rect 10538 3844 10590 4622
rect 10534 3840 10590 3844
rect 10694 3840 10696 4622
rect 10696 3840 10748 4622
rect 10748 3840 10750 4622
rect 10850 3844 10854 4622
rect 10854 3844 10906 4622
rect 10850 3840 10906 3844
rect 11010 3840 11012 4622
rect 11012 3840 11064 4622
rect 11064 3840 11066 4622
rect 11166 3844 11170 4622
rect 11170 3844 11222 4622
rect 11166 3840 11222 3844
rect 11326 3840 11328 4622
rect 11328 3840 11380 4622
rect 11380 3840 11382 4622
rect 11482 3844 11486 4622
rect 11486 3844 11538 4622
rect 11482 3840 11538 3844
rect 11642 3840 11644 4622
rect 11644 3840 11696 4622
rect 11696 3840 11698 4622
rect 11798 3844 11802 4622
rect 11802 3844 11854 4622
rect 11798 3840 11854 3844
rect 11958 3840 11960 4622
rect 11960 3840 12012 4622
rect 12012 3840 12014 4622
rect 12114 3844 12118 4622
rect 12118 3844 12170 4622
rect 12114 3840 12170 3844
rect 12274 3840 12276 4622
rect 12276 3840 12328 4622
rect 12328 3840 12330 4622
rect 12430 3844 12434 4622
rect 12434 3844 12486 4622
rect 12430 3840 12486 3844
rect 12590 3840 12592 4622
rect 12592 3840 12644 4622
rect 12644 3840 12646 4622
rect 12746 3844 12796 4622
rect 12796 3844 12802 4622
rect 12746 3840 12802 3844
rect 108 2934 110 3712
rect 110 2934 162 3712
rect 162 2934 164 3712
rect 266 2930 268 3712
rect 268 2930 320 3712
rect 320 2930 322 3712
rect 422 2932 426 3712
rect 426 2932 478 3712
rect 422 2930 478 2932
rect 582 2930 584 3712
rect 584 2930 636 3712
rect 636 2930 638 3712
rect 738 2932 742 3712
rect 742 2932 794 3712
rect 738 2930 794 2932
rect 898 2930 900 3712
rect 900 2930 952 3712
rect 952 2930 954 3712
rect 1054 2932 1058 3712
rect 1058 2932 1110 3712
rect 1054 2930 1110 2932
rect 1214 2930 1216 3712
rect 1216 2930 1268 3712
rect 1268 2930 1270 3712
rect 1370 2932 1374 3712
rect 1374 2932 1426 3712
rect 1370 2930 1426 2932
rect 1530 2930 1532 3712
rect 1532 2930 1584 3712
rect 1584 2930 1586 3712
rect 1686 2932 1690 3712
rect 1690 2932 1742 3712
rect 1686 2930 1742 2932
rect 1846 2930 1848 3712
rect 1848 2930 1900 3712
rect 1900 2930 1902 3712
rect 2002 2932 2006 3712
rect 2006 2932 2058 3712
rect 2002 2930 2058 2932
rect 2162 2930 2164 3712
rect 2164 2930 2216 3712
rect 2216 2930 2218 3712
rect 2318 2932 2322 3712
rect 2322 2932 2374 3712
rect 2318 2930 2374 2932
rect 2478 2930 2480 3712
rect 2480 2930 2532 3712
rect 2532 2930 2534 3712
rect 2634 2932 2638 3712
rect 2638 2932 2690 3712
rect 2634 2930 2690 2932
rect 2794 2930 2796 3712
rect 2796 2930 2848 3712
rect 2848 2930 2850 3712
rect 2950 2932 2954 3712
rect 2954 2932 3006 3712
rect 2950 2930 3006 2932
rect 3110 2930 3112 3712
rect 3112 2930 3164 3712
rect 3164 2930 3166 3712
rect 3266 2932 3270 3712
rect 3270 2932 3322 3712
rect 3266 2930 3322 2932
rect 3426 2930 3428 3712
rect 3428 2930 3480 3712
rect 3480 2930 3482 3712
rect 3582 2932 3586 3712
rect 3586 2932 3638 3712
rect 3582 2930 3638 2932
rect 3742 2930 3744 3712
rect 3744 2930 3796 3712
rect 3796 2930 3798 3712
rect 3898 2932 3902 3712
rect 3902 2932 3954 3712
rect 3898 2930 3954 2932
rect 4058 2930 4060 3712
rect 4060 2930 4112 3712
rect 4112 2930 4114 3712
rect 4214 2932 4218 3712
rect 4218 2932 4270 3712
rect 4214 2930 4270 2932
rect 4374 2930 4376 3712
rect 4376 2930 4428 3712
rect 4428 2930 4430 3712
rect 4530 2932 4534 3712
rect 4534 2932 4586 3712
rect 4530 2930 4586 2932
rect 4690 2930 4692 3712
rect 4692 2930 4744 3712
rect 4744 2930 4746 3712
rect 4846 2932 4850 3712
rect 4850 2932 4902 3712
rect 4846 2930 4902 2932
rect 5006 2930 5008 3712
rect 5008 2930 5060 3712
rect 5060 2930 5062 3712
rect 5162 2932 5166 3712
rect 5166 2932 5218 3712
rect 5162 2930 5218 2932
rect 5322 2930 5324 3712
rect 5324 2930 5376 3712
rect 5376 2930 5378 3712
rect 5478 2932 5482 3712
rect 5482 2932 5534 3712
rect 5478 2930 5534 2932
rect 5638 2930 5640 3712
rect 5640 2930 5692 3712
rect 5692 2930 5694 3712
rect 5794 2932 5798 3712
rect 5798 2932 5850 3712
rect 5794 2930 5850 2932
rect 5954 2930 5956 3712
rect 5956 2930 6008 3712
rect 6008 2930 6010 3712
rect 6110 2932 6114 3712
rect 6114 2932 6166 3712
rect 6110 2930 6166 2932
rect 6270 2930 6272 3712
rect 6272 2930 6324 3712
rect 6324 2930 6326 3712
rect 6426 2932 6430 3712
rect 6430 2932 6482 3712
rect 6426 2930 6482 2932
rect 6586 2930 6588 3712
rect 6588 2930 6640 3712
rect 6640 2930 6642 3712
rect 6742 2932 6746 3712
rect 6746 2932 6798 3712
rect 6742 2930 6798 2932
rect 6902 2930 6904 3712
rect 6904 2930 6956 3712
rect 6956 2930 6958 3712
rect 7058 2932 7062 3712
rect 7062 2932 7114 3712
rect 7058 2930 7114 2932
rect 7218 2930 7220 3712
rect 7220 2930 7272 3712
rect 7272 2930 7274 3712
rect 7374 2932 7378 3712
rect 7378 2932 7430 3712
rect 7374 2930 7430 2932
rect 7534 2930 7536 3712
rect 7536 2930 7588 3712
rect 7588 2930 7590 3712
rect 7690 2932 7694 3712
rect 7694 2932 7746 3712
rect 7690 2930 7746 2932
rect 7850 2930 7852 3712
rect 7852 2930 7904 3712
rect 7904 2930 7906 3712
rect 8006 2932 8010 3712
rect 8010 2932 8062 3712
rect 8006 2930 8062 2932
rect 8166 2930 8168 3712
rect 8168 2930 8220 3712
rect 8220 2930 8222 3712
rect 8322 2932 8326 3712
rect 8326 2932 8378 3712
rect 8322 2930 8378 2932
rect 8482 2930 8484 3712
rect 8484 2930 8536 3712
rect 8536 2930 8538 3712
rect 8638 2932 8642 3712
rect 8642 2932 8694 3712
rect 8638 2930 8694 2932
rect 8798 2930 8800 3712
rect 8800 2930 8852 3712
rect 8852 2930 8854 3712
rect 8954 2932 8958 3712
rect 8958 2932 9010 3712
rect 8954 2930 9010 2932
rect 9114 2930 9116 3712
rect 9116 2930 9168 3712
rect 9168 2930 9170 3712
rect 9270 2932 9274 3712
rect 9274 2932 9326 3712
rect 9270 2930 9326 2932
rect 9430 2930 9432 3712
rect 9432 2930 9484 3712
rect 9484 2930 9486 3712
rect 9586 2932 9590 3712
rect 9590 2932 9642 3712
rect 9586 2930 9642 2932
rect 9746 2930 9748 3712
rect 9748 2930 9800 3712
rect 9800 2930 9802 3712
rect 9902 2932 9906 3712
rect 9906 2932 9958 3712
rect 9902 2930 9958 2932
rect 10062 2930 10064 3712
rect 10064 2930 10116 3712
rect 10116 2930 10118 3712
rect 10218 2932 10222 3712
rect 10222 2932 10274 3712
rect 10218 2930 10274 2932
rect 10378 2930 10380 3712
rect 10380 2930 10432 3712
rect 10432 2930 10434 3712
rect 10534 2932 10538 3712
rect 10538 2932 10590 3712
rect 10534 2930 10590 2932
rect 10694 2930 10696 3712
rect 10696 2930 10748 3712
rect 10748 2930 10750 3712
rect 10850 2932 10854 3712
rect 10854 2932 10906 3712
rect 10850 2930 10906 2932
rect 11010 2930 11012 3712
rect 11012 2930 11064 3712
rect 11064 2930 11066 3712
rect 11166 2932 11170 3712
rect 11170 2932 11222 3712
rect 11166 2930 11222 2932
rect 11326 2930 11328 3712
rect 11328 2930 11380 3712
rect 11380 2930 11382 3712
rect 11482 2932 11486 3712
rect 11486 2932 11538 3712
rect 11482 2930 11538 2932
rect 11642 2930 11644 3712
rect 11644 2930 11696 3712
rect 11696 2930 11698 3712
rect 11798 2932 11802 3712
rect 11802 2932 11854 3712
rect 11798 2930 11854 2932
rect 11958 2930 11960 3712
rect 11960 2930 12012 3712
rect 12012 2930 12014 3712
rect 12114 2932 12118 3712
rect 12118 2932 12170 3712
rect 12114 2930 12170 2932
rect 12274 2930 12276 3712
rect 12276 2930 12328 3712
rect 12328 2930 12330 3712
rect 12430 2932 12434 3712
rect 12434 2932 12486 3712
rect 12430 2930 12486 2932
rect 12590 2930 12592 3712
rect 12592 2930 12644 3712
rect 12644 2930 12646 3712
rect 12746 2932 12796 3712
rect 12796 2932 12802 3712
rect 12746 2930 12802 2932
rect 108 2024 110 2802
rect 110 2024 162 2802
rect 162 2024 164 2802
rect 266 2020 268 2802
rect 268 2020 320 2802
rect 320 2020 322 2802
rect 422 2022 426 2802
rect 426 2022 478 2802
rect 422 2020 478 2022
rect 582 2020 584 2802
rect 584 2020 636 2802
rect 636 2020 638 2802
rect 738 2022 742 2802
rect 742 2022 794 2802
rect 738 2020 794 2022
rect 898 2020 900 2802
rect 900 2020 952 2802
rect 952 2020 954 2802
rect 1054 2022 1058 2802
rect 1058 2022 1110 2802
rect 1054 2020 1110 2022
rect 1214 2020 1216 2802
rect 1216 2020 1268 2802
rect 1268 2020 1270 2802
rect 1370 2022 1374 2802
rect 1374 2022 1426 2802
rect 1370 2020 1426 2022
rect 1530 2020 1532 2802
rect 1532 2020 1584 2802
rect 1584 2020 1586 2802
rect 1686 2022 1690 2802
rect 1690 2022 1742 2802
rect 1686 2020 1742 2022
rect 1846 2020 1848 2802
rect 1848 2020 1900 2802
rect 1900 2020 1902 2802
rect 2002 2022 2006 2802
rect 2006 2022 2058 2802
rect 2002 2020 2058 2022
rect 2162 2020 2164 2802
rect 2164 2020 2216 2802
rect 2216 2020 2218 2802
rect 2318 2022 2322 2802
rect 2322 2022 2374 2802
rect 2318 2020 2374 2022
rect 2478 2020 2480 2802
rect 2480 2020 2532 2802
rect 2532 2020 2534 2802
rect 2634 2022 2638 2802
rect 2638 2022 2690 2802
rect 2634 2020 2690 2022
rect 2794 2020 2796 2802
rect 2796 2020 2848 2802
rect 2848 2020 2850 2802
rect 2950 2022 2954 2802
rect 2954 2022 3006 2802
rect 2950 2020 3006 2022
rect 3110 2020 3112 2802
rect 3112 2020 3164 2802
rect 3164 2020 3166 2802
rect 3266 2022 3270 2802
rect 3270 2022 3322 2802
rect 3266 2020 3322 2022
rect 3426 2020 3428 2802
rect 3428 2020 3480 2802
rect 3480 2020 3482 2802
rect 3582 2022 3586 2802
rect 3586 2022 3638 2802
rect 3582 2020 3638 2022
rect 3742 2020 3744 2802
rect 3744 2020 3796 2802
rect 3796 2020 3798 2802
rect 3898 2022 3902 2802
rect 3902 2022 3954 2802
rect 3898 2020 3954 2022
rect 4058 2020 4060 2802
rect 4060 2020 4112 2802
rect 4112 2020 4114 2802
rect 4214 2022 4218 2802
rect 4218 2022 4270 2802
rect 4214 2020 4270 2022
rect 4374 2020 4376 2802
rect 4376 2020 4428 2802
rect 4428 2020 4430 2802
rect 4530 2022 4534 2802
rect 4534 2022 4586 2802
rect 4530 2020 4586 2022
rect 4690 2020 4692 2802
rect 4692 2020 4744 2802
rect 4744 2020 4746 2802
rect 4846 2022 4850 2802
rect 4850 2022 4902 2802
rect 4846 2020 4902 2022
rect 5006 2020 5008 2802
rect 5008 2020 5060 2802
rect 5060 2020 5062 2802
rect 5162 2022 5166 2802
rect 5166 2022 5218 2802
rect 5162 2020 5218 2022
rect 5322 2020 5324 2802
rect 5324 2020 5376 2802
rect 5376 2020 5378 2802
rect 5478 2022 5482 2802
rect 5482 2022 5534 2802
rect 5478 2020 5534 2022
rect 5638 2020 5640 2802
rect 5640 2020 5692 2802
rect 5692 2020 5694 2802
rect 5794 2022 5798 2802
rect 5798 2022 5850 2802
rect 5794 2020 5850 2022
rect 5954 2020 5956 2802
rect 5956 2020 6008 2802
rect 6008 2020 6010 2802
rect 6110 2022 6114 2802
rect 6114 2022 6166 2802
rect 6110 2020 6166 2022
rect 6270 2020 6272 2802
rect 6272 2020 6324 2802
rect 6324 2020 6326 2802
rect 6426 2022 6430 2802
rect 6430 2022 6482 2802
rect 6426 2020 6482 2022
rect 6586 2020 6588 2802
rect 6588 2020 6640 2802
rect 6640 2020 6642 2802
rect 6742 2022 6746 2802
rect 6746 2022 6798 2802
rect 6742 2020 6798 2022
rect 6902 2020 6904 2802
rect 6904 2020 6956 2802
rect 6956 2020 6958 2802
rect 7058 2022 7062 2802
rect 7062 2022 7114 2802
rect 7058 2020 7114 2022
rect 7218 2020 7220 2802
rect 7220 2020 7272 2802
rect 7272 2020 7274 2802
rect 7374 2022 7378 2802
rect 7378 2022 7430 2802
rect 7374 2020 7430 2022
rect 7534 2020 7536 2802
rect 7536 2020 7588 2802
rect 7588 2020 7590 2802
rect 7690 2022 7694 2802
rect 7694 2022 7746 2802
rect 7690 2020 7746 2022
rect 7850 2020 7852 2802
rect 7852 2020 7904 2802
rect 7904 2020 7906 2802
rect 8006 2022 8010 2802
rect 8010 2022 8062 2802
rect 8006 2020 8062 2022
rect 8166 2020 8168 2802
rect 8168 2020 8220 2802
rect 8220 2020 8222 2802
rect 8322 2022 8326 2802
rect 8326 2022 8378 2802
rect 8322 2020 8378 2022
rect 8482 2020 8484 2802
rect 8484 2020 8536 2802
rect 8536 2020 8538 2802
rect 8638 2022 8642 2802
rect 8642 2022 8694 2802
rect 8638 2020 8694 2022
rect 8798 2020 8800 2802
rect 8800 2020 8852 2802
rect 8852 2020 8854 2802
rect 8954 2022 8958 2802
rect 8958 2022 9010 2802
rect 8954 2020 9010 2022
rect 9114 2020 9116 2802
rect 9116 2020 9168 2802
rect 9168 2020 9170 2802
rect 9270 2022 9274 2802
rect 9274 2022 9326 2802
rect 9270 2020 9326 2022
rect 9430 2020 9432 2802
rect 9432 2020 9484 2802
rect 9484 2020 9486 2802
rect 9586 2022 9590 2802
rect 9590 2022 9642 2802
rect 9586 2020 9642 2022
rect 9746 2020 9748 2802
rect 9748 2020 9800 2802
rect 9800 2020 9802 2802
rect 9902 2022 9906 2802
rect 9906 2022 9958 2802
rect 9902 2020 9958 2022
rect 10062 2020 10064 2802
rect 10064 2020 10116 2802
rect 10116 2020 10118 2802
rect 10218 2022 10222 2802
rect 10222 2022 10274 2802
rect 10218 2020 10274 2022
rect 10378 2020 10380 2802
rect 10380 2020 10432 2802
rect 10432 2020 10434 2802
rect 10534 2022 10538 2802
rect 10538 2022 10590 2802
rect 10534 2020 10590 2022
rect 10694 2020 10696 2802
rect 10696 2020 10748 2802
rect 10748 2020 10750 2802
rect 10850 2022 10854 2802
rect 10854 2022 10906 2802
rect 10850 2020 10906 2022
rect 11010 2020 11012 2802
rect 11012 2020 11064 2802
rect 11064 2020 11066 2802
rect 11166 2022 11170 2802
rect 11170 2022 11222 2802
rect 11166 2020 11222 2022
rect 11326 2020 11328 2802
rect 11328 2020 11380 2802
rect 11380 2020 11382 2802
rect 11482 2022 11486 2802
rect 11486 2022 11538 2802
rect 11482 2020 11538 2022
rect 11642 2020 11644 2802
rect 11644 2020 11696 2802
rect 11696 2020 11698 2802
rect 11798 2022 11802 2802
rect 11802 2022 11854 2802
rect 11798 2020 11854 2022
rect 11958 2020 11960 2802
rect 11960 2020 12012 2802
rect 12012 2020 12014 2802
rect 12114 2022 12118 2802
rect 12118 2022 12170 2802
rect 12114 2020 12170 2022
rect 12274 2020 12276 2802
rect 12276 2020 12328 2802
rect 12328 2020 12330 2802
rect 12430 2022 12434 2802
rect 12434 2022 12486 2802
rect 12430 2020 12486 2022
rect 12590 2020 12592 2802
rect 12592 2020 12644 2802
rect 12644 2020 12646 2802
rect 12746 2022 12796 2802
rect 12796 2022 12802 2802
rect 12746 2020 12802 2022
rect 108 1114 110 1892
rect 110 1114 162 1892
rect 162 1114 164 1892
rect 266 1110 268 1892
rect 268 1110 320 1892
rect 320 1110 322 1892
rect 422 1112 426 1892
rect 426 1112 478 1892
rect 422 1110 478 1112
rect 582 1110 584 1892
rect 584 1110 636 1892
rect 636 1110 638 1892
rect 738 1112 742 1892
rect 742 1112 794 1892
rect 738 1110 794 1112
rect 898 1110 900 1892
rect 900 1110 952 1892
rect 952 1110 954 1892
rect 1054 1112 1058 1892
rect 1058 1112 1110 1892
rect 1054 1110 1110 1112
rect 1214 1110 1216 1892
rect 1216 1110 1268 1892
rect 1268 1110 1270 1892
rect 1370 1112 1374 1892
rect 1374 1112 1426 1892
rect 1370 1110 1426 1112
rect 1530 1110 1532 1892
rect 1532 1110 1584 1892
rect 1584 1110 1586 1892
rect 1686 1112 1690 1892
rect 1690 1112 1742 1892
rect 1686 1110 1742 1112
rect 1846 1110 1848 1892
rect 1848 1110 1900 1892
rect 1900 1110 1902 1892
rect 2002 1112 2006 1892
rect 2006 1112 2058 1892
rect 2002 1110 2058 1112
rect 2162 1110 2164 1892
rect 2164 1110 2216 1892
rect 2216 1110 2218 1892
rect 2318 1112 2322 1892
rect 2322 1112 2374 1892
rect 2318 1110 2374 1112
rect 2478 1110 2480 1892
rect 2480 1110 2532 1892
rect 2532 1110 2534 1892
rect 2634 1112 2638 1892
rect 2638 1112 2690 1892
rect 2634 1110 2690 1112
rect 2794 1110 2796 1892
rect 2796 1110 2848 1892
rect 2848 1110 2850 1892
rect 2950 1112 2954 1892
rect 2954 1112 3006 1892
rect 2950 1110 3006 1112
rect 3110 1110 3112 1892
rect 3112 1110 3164 1892
rect 3164 1110 3166 1892
rect 3266 1112 3270 1892
rect 3270 1112 3322 1892
rect 3266 1110 3322 1112
rect 3426 1110 3428 1892
rect 3428 1110 3480 1892
rect 3480 1110 3482 1892
rect 3582 1112 3586 1892
rect 3586 1112 3638 1892
rect 3582 1110 3638 1112
rect 3742 1110 3744 1892
rect 3744 1110 3796 1892
rect 3796 1110 3798 1892
rect 3898 1112 3902 1892
rect 3902 1112 3954 1892
rect 3898 1110 3954 1112
rect 4058 1110 4060 1892
rect 4060 1110 4112 1892
rect 4112 1110 4114 1892
rect 4214 1112 4218 1892
rect 4218 1112 4270 1892
rect 4214 1110 4270 1112
rect 4374 1110 4376 1892
rect 4376 1110 4428 1892
rect 4428 1110 4430 1892
rect 4530 1112 4534 1892
rect 4534 1112 4586 1892
rect 4530 1110 4586 1112
rect 4690 1110 4692 1892
rect 4692 1110 4744 1892
rect 4744 1110 4746 1892
rect 4846 1112 4850 1892
rect 4850 1112 4902 1892
rect 4846 1110 4902 1112
rect 5006 1110 5008 1892
rect 5008 1110 5060 1892
rect 5060 1110 5062 1892
rect 5162 1112 5166 1892
rect 5166 1112 5218 1892
rect 5162 1110 5218 1112
rect 5322 1110 5324 1892
rect 5324 1110 5376 1892
rect 5376 1110 5378 1892
rect 5478 1112 5482 1892
rect 5482 1112 5534 1892
rect 5478 1110 5534 1112
rect 5638 1110 5640 1892
rect 5640 1110 5692 1892
rect 5692 1110 5694 1892
rect 5794 1112 5798 1892
rect 5798 1112 5850 1892
rect 5794 1110 5850 1112
rect 5954 1110 5956 1892
rect 5956 1110 6008 1892
rect 6008 1110 6010 1892
rect 6110 1112 6114 1892
rect 6114 1112 6166 1892
rect 6110 1110 6166 1112
rect 6270 1110 6272 1892
rect 6272 1110 6324 1892
rect 6324 1110 6326 1892
rect 6426 1112 6430 1892
rect 6430 1112 6482 1892
rect 6426 1110 6482 1112
rect 6586 1110 6588 1892
rect 6588 1110 6640 1892
rect 6640 1110 6642 1892
rect 6742 1112 6746 1892
rect 6746 1112 6798 1892
rect 6742 1110 6798 1112
rect 6902 1110 6904 1892
rect 6904 1110 6956 1892
rect 6956 1110 6958 1892
rect 7058 1112 7062 1892
rect 7062 1112 7114 1892
rect 7058 1110 7114 1112
rect 7218 1110 7220 1892
rect 7220 1110 7272 1892
rect 7272 1110 7274 1892
rect 7374 1112 7378 1892
rect 7378 1112 7430 1892
rect 7374 1110 7430 1112
rect 7534 1110 7536 1892
rect 7536 1110 7588 1892
rect 7588 1110 7590 1892
rect 7690 1112 7694 1892
rect 7694 1112 7746 1892
rect 7690 1110 7746 1112
rect 7850 1110 7852 1892
rect 7852 1110 7904 1892
rect 7904 1110 7906 1892
rect 8006 1112 8010 1892
rect 8010 1112 8062 1892
rect 8006 1110 8062 1112
rect 8166 1110 8168 1892
rect 8168 1110 8220 1892
rect 8220 1110 8222 1892
rect 8322 1112 8326 1892
rect 8326 1112 8378 1892
rect 8322 1110 8378 1112
rect 8482 1110 8484 1892
rect 8484 1110 8536 1892
rect 8536 1110 8538 1892
rect 8638 1112 8642 1892
rect 8642 1112 8694 1892
rect 8638 1110 8694 1112
rect 8798 1110 8800 1892
rect 8800 1110 8852 1892
rect 8852 1110 8854 1892
rect 8954 1112 8958 1892
rect 8958 1112 9010 1892
rect 8954 1110 9010 1112
rect 9114 1110 9116 1892
rect 9116 1110 9168 1892
rect 9168 1110 9170 1892
rect 9270 1112 9274 1892
rect 9274 1112 9326 1892
rect 9270 1110 9326 1112
rect 9430 1110 9432 1892
rect 9432 1110 9484 1892
rect 9484 1110 9486 1892
rect 9586 1112 9590 1892
rect 9590 1112 9642 1892
rect 9586 1110 9642 1112
rect 9746 1110 9748 1892
rect 9748 1110 9800 1892
rect 9800 1110 9802 1892
rect 9902 1112 9906 1892
rect 9906 1112 9958 1892
rect 9902 1110 9958 1112
rect 10062 1110 10064 1892
rect 10064 1110 10116 1892
rect 10116 1110 10118 1892
rect 10218 1112 10222 1892
rect 10222 1112 10274 1892
rect 10218 1110 10274 1112
rect 10378 1110 10380 1892
rect 10380 1110 10432 1892
rect 10432 1110 10434 1892
rect 10534 1112 10538 1892
rect 10538 1112 10590 1892
rect 10534 1110 10590 1112
rect 10694 1110 10696 1892
rect 10696 1110 10748 1892
rect 10748 1110 10750 1892
rect 10850 1112 10854 1892
rect 10854 1112 10906 1892
rect 10850 1110 10906 1112
rect 11010 1110 11012 1892
rect 11012 1110 11064 1892
rect 11064 1110 11066 1892
rect 11166 1112 11170 1892
rect 11170 1112 11222 1892
rect 11166 1110 11222 1112
rect 11326 1110 11328 1892
rect 11328 1110 11380 1892
rect 11380 1110 11382 1892
rect 11482 1112 11486 1892
rect 11486 1112 11538 1892
rect 11482 1110 11538 1112
rect 11642 1110 11644 1892
rect 11644 1110 11696 1892
rect 11696 1110 11698 1892
rect 11798 1112 11802 1892
rect 11802 1112 11854 1892
rect 11798 1110 11854 1112
rect 11958 1110 11960 1892
rect 11960 1110 12012 1892
rect 12012 1110 12014 1892
rect 12114 1112 12118 1892
rect 12118 1112 12170 1892
rect 12114 1110 12170 1112
rect 12274 1110 12276 1892
rect 12276 1110 12328 1892
rect 12328 1110 12330 1892
rect 12430 1112 12434 1892
rect 12434 1112 12486 1892
rect 12430 1110 12486 1112
rect 12590 1110 12592 1892
rect 12592 1110 12644 1892
rect 12644 1110 12646 1892
rect 12746 1112 12796 1892
rect 12796 1112 12802 1892
rect 12746 1110 12802 1112
rect 108 204 110 982
rect 110 204 162 982
rect 162 204 164 982
rect 266 980 322 982
rect 266 202 268 980
rect 268 202 320 980
rect 320 202 322 980
rect 266 200 322 202
rect 422 202 426 982
rect 426 202 478 982
rect 422 200 478 202
rect 582 980 638 982
rect 582 202 584 980
rect 584 202 636 980
rect 636 202 638 980
rect 582 200 638 202
rect 738 202 742 982
rect 742 202 794 982
rect 738 200 794 202
rect 898 980 954 982
rect 898 202 900 980
rect 900 202 952 980
rect 952 202 954 980
rect 898 200 954 202
rect 1054 202 1058 982
rect 1058 202 1110 982
rect 1054 200 1110 202
rect 1214 980 1270 982
rect 1214 202 1216 980
rect 1216 202 1268 980
rect 1268 202 1270 980
rect 1214 200 1270 202
rect 1370 202 1374 982
rect 1374 202 1426 982
rect 1370 200 1426 202
rect 1530 980 1586 982
rect 1530 202 1532 980
rect 1532 202 1584 980
rect 1584 202 1586 980
rect 1530 200 1586 202
rect 1686 202 1690 982
rect 1690 202 1742 982
rect 1686 200 1742 202
rect 1846 980 1902 982
rect 1846 202 1848 980
rect 1848 202 1900 980
rect 1900 202 1902 980
rect 1846 200 1902 202
rect 2002 202 2006 982
rect 2006 202 2058 982
rect 2002 200 2058 202
rect 2162 980 2218 982
rect 2162 202 2164 980
rect 2164 202 2216 980
rect 2216 202 2218 980
rect 2162 200 2218 202
rect 2318 202 2322 982
rect 2322 202 2374 982
rect 2318 200 2374 202
rect 2478 980 2534 982
rect 2478 202 2480 980
rect 2480 202 2532 980
rect 2532 202 2534 980
rect 2478 200 2534 202
rect 2634 202 2638 982
rect 2638 202 2690 982
rect 2634 200 2690 202
rect 2794 980 2850 982
rect 2794 202 2796 980
rect 2796 202 2848 980
rect 2848 202 2850 980
rect 2794 200 2850 202
rect 2950 202 2954 982
rect 2954 202 3006 982
rect 2950 200 3006 202
rect 3110 980 3166 982
rect 3110 202 3112 980
rect 3112 202 3164 980
rect 3164 202 3166 980
rect 3110 200 3166 202
rect 3266 202 3270 982
rect 3270 202 3322 982
rect 3266 200 3322 202
rect 3426 980 3482 982
rect 3426 202 3428 980
rect 3428 202 3480 980
rect 3480 202 3482 980
rect 3426 200 3482 202
rect 3582 202 3586 982
rect 3586 202 3638 982
rect 3582 200 3638 202
rect 3742 980 3798 982
rect 3742 202 3744 980
rect 3744 202 3796 980
rect 3796 202 3798 980
rect 3742 200 3798 202
rect 3898 202 3902 982
rect 3902 202 3954 982
rect 3898 200 3954 202
rect 4058 980 4114 982
rect 4058 202 4060 980
rect 4060 202 4112 980
rect 4112 202 4114 980
rect 4058 200 4114 202
rect 4214 202 4218 982
rect 4218 202 4270 982
rect 4214 200 4270 202
rect 4374 980 4430 982
rect 4374 202 4376 980
rect 4376 202 4428 980
rect 4428 202 4430 980
rect 4374 200 4430 202
rect 4530 202 4534 982
rect 4534 202 4586 982
rect 4530 200 4586 202
rect 4690 980 4746 982
rect 4690 202 4692 980
rect 4692 202 4744 980
rect 4744 202 4746 980
rect 4690 200 4746 202
rect 4846 202 4850 982
rect 4850 202 4902 982
rect 4846 200 4902 202
rect 5006 980 5062 982
rect 5006 202 5008 980
rect 5008 202 5060 980
rect 5060 202 5062 980
rect 5006 200 5062 202
rect 5162 202 5166 982
rect 5166 202 5218 982
rect 5162 200 5218 202
rect 5322 980 5378 982
rect 5322 202 5324 980
rect 5324 202 5376 980
rect 5376 202 5378 980
rect 5322 200 5378 202
rect 5478 202 5482 982
rect 5482 202 5534 982
rect 5478 200 5534 202
rect 5638 980 5694 982
rect 5638 202 5640 980
rect 5640 202 5692 980
rect 5692 202 5694 980
rect 5638 200 5694 202
rect 5794 202 5798 982
rect 5798 202 5850 982
rect 5794 200 5850 202
rect 5954 980 6010 982
rect 5954 202 5956 980
rect 5956 202 6008 980
rect 6008 202 6010 980
rect 5954 200 6010 202
rect 6110 202 6114 982
rect 6114 202 6166 982
rect 6110 200 6166 202
rect 6270 980 6326 982
rect 6270 202 6272 980
rect 6272 202 6324 980
rect 6324 202 6326 980
rect 6270 200 6326 202
rect 6426 202 6430 982
rect 6430 202 6482 982
rect 6426 200 6482 202
rect 6586 980 6642 982
rect 6586 202 6588 980
rect 6588 202 6640 980
rect 6640 202 6642 980
rect 6586 200 6642 202
rect 6742 202 6746 982
rect 6746 202 6798 982
rect 6742 200 6798 202
rect 6902 980 6958 982
rect 6902 202 6904 980
rect 6904 202 6956 980
rect 6956 202 6958 980
rect 6902 200 6958 202
rect 7058 202 7062 982
rect 7062 202 7114 982
rect 7058 200 7114 202
rect 7218 980 7274 982
rect 7218 202 7220 980
rect 7220 202 7272 980
rect 7272 202 7274 980
rect 7218 200 7274 202
rect 7374 202 7378 982
rect 7378 202 7430 982
rect 7374 200 7430 202
rect 7534 980 7590 982
rect 7534 202 7536 980
rect 7536 202 7588 980
rect 7588 202 7590 980
rect 7534 200 7590 202
rect 7690 202 7694 982
rect 7694 202 7746 982
rect 7690 200 7746 202
rect 7850 980 7906 982
rect 7850 202 7852 980
rect 7852 202 7904 980
rect 7904 202 7906 980
rect 7850 200 7906 202
rect 8006 202 8010 982
rect 8010 202 8062 982
rect 8006 200 8062 202
rect 8166 980 8222 982
rect 8166 202 8168 980
rect 8168 202 8220 980
rect 8220 202 8222 980
rect 8166 200 8222 202
rect 8322 202 8326 982
rect 8326 202 8378 982
rect 8322 200 8378 202
rect 8482 980 8538 982
rect 8482 202 8484 980
rect 8484 202 8536 980
rect 8536 202 8538 980
rect 8482 200 8538 202
rect 8638 202 8642 982
rect 8642 202 8694 982
rect 8638 200 8694 202
rect 8798 980 8854 982
rect 8798 202 8800 980
rect 8800 202 8852 980
rect 8852 202 8854 980
rect 8798 200 8854 202
rect 8954 202 8958 982
rect 8958 202 9010 982
rect 8954 200 9010 202
rect 9114 980 9170 982
rect 9114 202 9116 980
rect 9116 202 9168 980
rect 9168 202 9170 980
rect 9114 200 9170 202
rect 9270 202 9274 982
rect 9274 202 9326 982
rect 9270 200 9326 202
rect 9430 980 9486 982
rect 9430 202 9432 980
rect 9432 202 9484 980
rect 9484 202 9486 980
rect 9430 200 9486 202
rect 9586 202 9590 982
rect 9590 202 9642 982
rect 9586 200 9642 202
rect 9746 980 9802 982
rect 9746 202 9748 980
rect 9748 202 9800 980
rect 9800 202 9802 980
rect 9746 200 9802 202
rect 9902 202 9906 982
rect 9906 202 9958 982
rect 9902 200 9958 202
rect 10062 980 10118 982
rect 10062 202 10064 980
rect 10064 202 10116 980
rect 10116 202 10118 980
rect 10062 200 10118 202
rect 10218 202 10222 982
rect 10222 202 10274 982
rect 10218 200 10274 202
rect 10378 980 10434 982
rect 10378 202 10380 980
rect 10380 202 10432 980
rect 10432 202 10434 980
rect 10378 200 10434 202
rect 10534 202 10538 982
rect 10538 202 10590 982
rect 10534 200 10590 202
rect 10694 980 10750 982
rect 10694 202 10696 980
rect 10696 202 10748 980
rect 10748 202 10750 980
rect 10694 200 10750 202
rect 10850 202 10854 982
rect 10854 202 10906 982
rect 10850 200 10906 202
rect 11010 980 11066 982
rect 11010 202 11012 980
rect 11012 202 11064 980
rect 11064 202 11066 980
rect 11010 200 11066 202
rect 11166 202 11170 982
rect 11170 202 11222 982
rect 11166 200 11222 202
rect 11326 980 11382 982
rect 11326 202 11328 980
rect 11328 202 11380 980
rect 11380 202 11382 980
rect 11326 200 11382 202
rect 11482 202 11486 982
rect 11486 202 11538 982
rect 11482 200 11538 202
rect 11642 980 11698 982
rect 11642 202 11644 980
rect 11644 202 11696 980
rect 11696 202 11698 980
rect 11642 200 11698 202
rect 11798 202 11802 982
rect 11802 202 11854 982
rect 11798 200 11854 202
rect 11958 980 12014 982
rect 11958 202 11960 980
rect 11960 202 12012 980
rect 12012 202 12014 980
rect 11958 200 12014 202
rect 12114 202 12118 982
rect 12118 202 12170 982
rect 12114 200 12170 202
rect 12274 980 12330 982
rect 12274 202 12276 980
rect 12276 202 12328 980
rect 12328 202 12330 980
rect 12274 200 12330 202
rect 12430 202 12434 982
rect 12434 202 12486 982
rect 12430 200 12486 202
rect 12590 980 12646 982
rect 12590 202 12592 980
rect 12592 202 12644 980
rect 12644 202 12646 980
rect 12590 200 12646 202
rect 12746 202 12796 982
rect 12796 202 12802 982
rect 12746 200 12802 202
<< metal3 >>
rect 102 4632 166 4890
rect 260 4632 324 4890
rect 418 4632 482 4890
rect 576 4632 640 4890
rect 734 4632 798 4890
rect 892 4632 956 4890
rect 1050 4632 1114 4890
rect 1208 4632 1272 4890
rect 1366 4632 1430 4890
rect 1524 4632 1588 4890
rect 1682 4632 1746 4890
rect 1840 4632 1904 4890
rect 1998 4632 2062 4890
rect 2156 4632 2220 4890
rect 2314 4632 2378 4890
rect 2472 4632 2536 4890
rect 2630 4632 2694 4890
rect 2788 4632 2852 4890
rect 2946 4632 3010 4890
rect 3104 4632 3168 4890
rect 3262 4632 3326 4890
rect 3420 4632 3484 4890
rect 3578 4632 3642 4890
rect 3736 4632 3800 4890
rect 3894 4632 3958 4890
rect 4052 4632 4116 4890
rect 4210 4632 4274 4890
rect 4368 4632 4432 4890
rect 4526 4632 4590 4890
rect 4684 4632 4748 4890
rect 4842 4632 4906 4890
rect 5000 4632 5064 4890
rect 5158 4632 5222 4890
rect 5316 4632 5380 4890
rect 5474 4632 5538 4890
rect 5632 4632 5696 4890
rect 5790 4632 5854 4890
rect 5948 4632 6012 4890
rect 6106 4632 6170 4890
rect 6264 4632 6328 4890
rect 6422 4632 6486 4890
rect 6580 4632 6644 4890
rect 6738 4632 6802 4890
rect 6896 4632 6960 4890
rect 7054 4632 7118 4890
rect 7212 4632 7276 4890
rect 7370 4632 7434 4890
rect 7528 4632 7592 4890
rect 7686 4632 7750 4890
rect 7844 4632 7908 4890
rect 8002 4632 8066 4890
rect 8160 4632 8224 4890
rect 8318 4632 8382 4890
rect 8476 4632 8540 4890
rect 8634 4632 8698 4890
rect 8792 4632 8856 4890
rect 8950 4632 9014 4890
rect 9108 4632 9172 4890
rect 9266 4632 9330 4890
rect 9424 4632 9488 4890
rect 9582 4632 9646 4890
rect 9740 4632 9804 4890
rect 9898 4632 9962 4890
rect 10056 4632 10120 4890
rect 10214 4632 10278 4890
rect 10372 4632 10436 4890
rect 10530 4632 10594 4890
rect 10688 4632 10752 4890
rect 10846 4632 10910 4890
rect 11004 4632 11068 4890
rect 11162 4632 11226 4890
rect 11320 4632 11384 4890
rect 11478 4632 11542 4890
rect 11636 4632 11700 4890
rect 11794 4632 11858 4890
rect 11952 4632 12016 4890
rect 12110 4632 12174 4890
rect 12268 4632 12332 4890
rect 12426 4632 12490 4890
rect 12584 4632 12648 4890
rect 12742 4632 12806 4890
rect 98 4622 172 4632
rect 98 3844 108 4622
rect 164 3844 172 4622
rect 98 3834 172 3844
rect 256 4622 328 4632
rect 256 3840 266 4622
rect 322 3840 328 4622
rect 102 3722 166 3834
rect 256 3830 328 3840
rect 412 4622 488 4632
rect 412 3840 422 4622
rect 478 3840 488 4622
rect 412 3830 488 3840
rect 572 4622 644 4632
rect 572 3840 582 4622
rect 638 3840 644 4622
rect 572 3830 644 3840
rect 728 4622 804 4632
rect 728 3840 738 4622
rect 794 3840 804 4622
rect 728 3830 804 3840
rect 888 4622 960 4632
rect 888 3840 898 4622
rect 954 3840 960 4622
rect 888 3830 960 3840
rect 1044 4622 1120 4632
rect 1044 3840 1054 4622
rect 1110 3840 1120 4622
rect 1044 3830 1120 3840
rect 1204 4622 1276 4632
rect 1204 3840 1214 4622
rect 1270 3840 1276 4622
rect 1204 3830 1276 3840
rect 1360 4622 1436 4632
rect 1360 3840 1370 4622
rect 1426 3840 1436 4622
rect 1360 3830 1436 3840
rect 1520 4622 1592 4632
rect 1520 3840 1530 4622
rect 1586 3840 1592 4622
rect 1520 3830 1592 3840
rect 1676 4622 1752 4632
rect 1676 3840 1686 4622
rect 1742 3840 1752 4622
rect 1676 3830 1752 3840
rect 1836 4622 1908 4632
rect 1836 3840 1846 4622
rect 1902 3840 1908 4622
rect 1836 3830 1908 3840
rect 1992 4622 2068 4632
rect 1992 3840 2002 4622
rect 2058 3840 2068 4622
rect 1992 3830 2068 3840
rect 2152 4622 2224 4632
rect 2152 3840 2162 4622
rect 2218 3840 2224 4622
rect 2152 3830 2224 3840
rect 2308 4622 2384 4632
rect 2308 3840 2318 4622
rect 2374 3840 2384 4622
rect 2308 3830 2384 3840
rect 2468 4622 2540 4632
rect 2468 3840 2478 4622
rect 2534 3840 2540 4622
rect 2468 3830 2540 3840
rect 2624 4622 2700 4632
rect 2624 3840 2634 4622
rect 2690 3840 2700 4622
rect 2624 3830 2700 3840
rect 2784 4622 2856 4632
rect 2784 3840 2794 4622
rect 2850 3840 2856 4622
rect 2784 3830 2856 3840
rect 2940 4622 3016 4632
rect 2940 3840 2950 4622
rect 3006 3840 3016 4622
rect 2940 3830 3016 3840
rect 3100 4622 3172 4632
rect 3100 3840 3110 4622
rect 3166 3840 3172 4622
rect 3100 3830 3172 3840
rect 3256 4622 3332 4632
rect 3256 3840 3266 4622
rect 3322 3840 3332 4622
rect 3256 3830 3332 3840
rect 3416 4622 3488 4632
rect 3416 3840 3426 4622
rect 3482 3840 3488 4622
rect 3416 3830 3488 3840
rect 3572 4622 3648 4632
rect 3572 3840 3582 4622
rect 3638 3840 3648 4622
rect 3572 3830 3648 3840
rect 3732 4622 3804 4632
rect 3732 3840 3742 4622
rect 3798 3840 3804 4622
rect 3732 3830 3804 3840
rect 3888 4622 3964 4632
rect 3888 3840 3898 4622
rect 3954 3840 3964 4622
rect 3888 3830 3964 3840
rect 4048 4622 4120 4632
rect 4048 3840 4058 4622
rect 4114 3840 4120 4622
rect 4048 3830 4120 3840
rect 4204 4622 4280 4632
rect 4204 3840 4214 4622
rect 4270 3840 4280 4622
rect 4204 3830 4280 3840
rect 4364 4622 4436 4632
rect 4364 3840 4374 4622
rect 4430 3840 4436 4622
rect 4364 3830 4436 3840
rect 4520 4622 4596 4632
rect 4520 3840 4530 4622
rect 4586 3840 4596 4622
rect 4520 3830 4596 3840
rect 4680 4622 4752 4632
rect 4680 3840 4690 4622
rect 4746 3840 4752 4622
rect 4680 3830 4752 3840
rect 4836 4622 4912 4632
rect 4836 3840 4846 4622
rect 4902 3840 4912 4622
rect 4836 3830 4912 3840
rect 4996 4622 5068 4632
rect 4996 3840 5006 4622
rect 5062 3840 5068 4622
rect 4996 3830 5068 3840
rect 5152 4622 5228 4632
rect 5152 3840 5162 4622
rect 5218 3840 5228 4622
rect 5152 3830 5228 3840
rect 5312 4622 5384 4632
rect 5312 3840 5322 4622
rect 5378 3840 5384 4622
rect 5312 3830 5384 3840
rect 5468 4622 5544 4632
rect 5468 3840 5478 4622
rect 5534 3840 5544 4622
rect 5468 3830 5544 3840
rect 5628 4622 5700 4632
rect 5628 3840 5638 4622
rect 5694 3840 5700 4622
rect 5628 3830 5700 3840
rect 5784 4622 5860 4632
rect 5784 3840 5794 4622
rect 5850 3840 5860 4622
rect 5784 3830 5860 3840
rect 5944 4622 6016 4632
rect 5944 3840 5954 4622
rect 6010 3840 6016 4622
rect 5944 3830 6016 3840
rect 6100 4622 6176 4632
rect 6100 3840 6110 4622
rect 6166 3840 6176 4622
rect 6100 3830 6176 3840
rect 6260 4622 6332 4632
rect 6260 3840 6270 4622
rect 6326 3840 6332 4622
rect 6260 3830 6332 3840
rect 6416 4622 6492 4632
rect 6416 3840 6426 4622
rect 6482 3840 6492 4622
rect 6416 3830 6492 3840
rect 6576 4622 6648 4632
rect 6576 3840 6586 4622
rect 6642 3840 6648 4622
rect 6576 3830 6648 3840
rect 6732 4622 6808 4632
rect 6732 3840 6742 4622
rect 6798 3840 6808 4622
rect 6732 3830 6808 3840
rect 6892 4622 6964 4632
rect 6892 3840 6902 4622
rect 6958 3840 6964 4622
rect 6892 3830 6964 3840
rect 7048 4622 7124 4632
rect 7048 3840 7058 4622
rect 7114 3840 7124 4622
rect 7048 3830 7124 3840
rect 7208 4622 7280 4632
rect 7208 3840 7218 4622
rect 7274 3840 7280 4622
rect 7208 3830 7280 3840
rect 7364 4622 7440 4632
rect 7364 3840 7374 4622
rect 7430 3840 7440 4622
rect 7364 3830 7440 3840
rect 7524 4622 7596 4632
rect 7524 3840 7534 4622
rect 7590 3840 7596 4622
rect 7524 3830 7596 3840
rect 7680 4622 7756 4632
rect 7680 3840 7690 4622
rect 7746 3840 7756 4622
rect 7680 3830 7756 3840
rect 7840 4622 7912 4632
rect 7840 3840 7850 4622
rect 7906 3840 7912 4622
rect 7840 3830 7912 3840
rect 7996 4622 8072 4632
rect 7996 3840 8006 4622
rect 8062 3840 8072 4622
rect 7996 3830 8072 3840
rect 8156 4622 8228 4632
rect 8156 3840 8166 4622
rect 8222 3840 8228 4622
rect 8156 3830 8228 3840
rect 8312 4622 8388 4632
rect 8312 3840 8322 4622
rect 8378 3840 8388 4622
rect 8312 3830 8388 3840
rect 8472 4622 8544 4632
rect 8472 3840 8482 4622
rect 8538 3840 8544 4622
rect 8472 3830 8544 3840
rect 8628 4622 8704 4632
rect 8628 3840 8638 4622
rect 8694 3840 8704 4622
rect 8628 3830 8704 3840
rect 8788 4622 8860 4632
rect 8788 3840 8798 4622
rect 8854 3840 8860 4622
rect 8788 3830 8860 3840
rect 8944 4622 9020 4632
rect 8944 3840 8954 4622
rect 9010 3840 9020 4622
rect 8944 3830 9020 3840
rect 9104 4622 9176 4632
rect 9104 3840 9114 4622
rect 9170 3840 9176 4622
rect 9104 3830 9176 3840
rect 9260 4622 9336 4632
rect 9260 3840 9270 4622
rect 9326 3840 9336 4622
rect 9260 3830 9336 3840
rect 9420 4622 9492 4632
rect 9420 3840 9430 4622
rect 9486 3840 9492 4622
rect 9420 3830 9492 3840
rect 9576 4622 9652 4632
rect 9576 3840 9586 4622
rect 9642 3840 9652 4622
rect 9576 3830 9652 3840
rect 9736 4622 9808 4632
rect 9736 3840 9746 4622
rect 9802 3840 9808 4622
rect 9736 3830 9808 3840
rect 9892 4622 9968 4632
rect 9892 3840 9902 4622
rect 9958 3840 9968 4622
rect 9892 3830 9968 3840
rect 10052 4622 10124 4632
rect 10052 3840 10062 4622
rect 10118 3840 10124 4622
rect 10052 3830 10124 3840
rect 10208 4622 10284 4632
rect 10208 3840 10218 4622
rect 10274 3840 10284 4622
rect 10208 3830 10284 3840
rect 10368 4622 10440 4632
rect 10368 3840 10378 4622
rect 10434 3840 10440 4622
rect 10368 3830 10440 3840
rect 10524 4622 10600 4632
rect 10524 3840 10534 4622
rect 10590 3840 10600 4622
rect 10524 3830 10600 3840
rect 10684 4622 10756 4632
rect 10684 3840 10694 4622
rect 10750 3840 10756 4622
rect 10684 3830 10756 3840
rect 10840 4622 10916 4632
rect 10840 3840 10850 4622
rect 10906 3840 10916 4622
rect 10840 3830 10916 3840
rect 11000 4622 11072 4632
rect 11000 3840 11010 4622
rect 11066 3840 11072 4622
rect 11000 3830 11072 3840
rect 11156 4622 11232 4632
rect 11156 3840 11166 4622
rect 11222 3840 11232 4622
rect 11156 3830 11232 3840
rect 11316 4622 11388 4632
rect 11316 3840 11326 4622
rect 11382 3840 11388 4622
rect 11316 3830 11388 3840
rect 11472 4622 11548 4632
rect 11472 3840 11482 4622
rect 11538 3840 11548 4622
rect 11472 3830 11548 3840
rect 11632 4622 11704 4632
rect 11632 3840 11642 4622
rect 11698 3840 11704 4622
rect 11632 3830 11704 3840
rect 11788 4622 11864 4632
rect 11788 3840 11798 4622
rect 11854 3840 11864 4622
rect 11788 3830 11864 3840
rect 11948 4622 12020 4632
rect 11948 3840 11958 4622
rect 12014 3840 12020 4622
rect 11948 3830 12020 3840
rect 12104 4622 12180 4632
rect 12104 3840 12114 4622
rect 12170 3840 12180 4622
rect 12104 3830 12180 3840
rect 12264 4622 12336 4632
rect 12264 3840 12274 4622
rect 12330 3840 12336 4622
rect 12264 3830 12336 3840
rect 12420 4622 12496 4632
rect 12420 3840 12430 4622
rect 12486 3840 12496 4622
rect 12420 3830 12496 3840
rect 12580 4622 12652 4632
rect 12580 3840 12590 4622
rect 12646 3840 12652 4622
rect 12580 3830 12652 3840
rect 12736 4622 12812 4632
rect 12736 3840 12746 4622
rect 12802 3840 12812 4622
rect 12736 3830 12812 3840
rect 260 3722 324 3830
rect 418 3722 482 3830
rect 576 3722 640 3830
rect 734 3722 798 3830
rect 892 3722 956 3830
rect 1050 3722 1114 3830
rect 1208 3722 1272 3830
rect 1366 3722 1430 3830
rect 1524 3722 1588 3830
rect 1682 3722 1746 3830
rect 1840 3722 1904 3830
rect 1998 3722 2062 3830
rect 2156 3722 2220 3830
rect 2314 3722 2378 3830
rect 2472 3722 2536 3830
rect 2630 3722 2694 3830
rect 2788 3722 2852 3830
rect 2946 3722 3010 3830
rect 3104 3722 3168 3830
rect 3262 3722 3326 3830
rect 3420 3722 3484 3830
rect 3578 3722 3642 3830
rect 3736 3722 3800 3830
rect 3894 3722 3958 3830
rect 4052 3722 4116 3830
rect 4210 3722 4274 3830
rect 4368 3722 4432 3830
rect 4526 3722 4590 3830
rect 4684 3722 4748 3830
rect 4842 3722 4906 3830
rect 5000 3722 5064 3830
rect 5158 3722 5222 3830
rect 5316 3722 5380 3830
rect 5474 3722 5538 3830
rect 5632 3722 5696 3830
rect 5790 3722 5854 3830
rect 5948 3722 6012 3830
rect 6106 3722 6170 3830
rect 6264 3722 6328 3830
rect 6422 3722 6486 3830
rect 6580 3722 6644 3830
rect 6738 3722 6802 3830
rect 6896 3722 6960 3830
rect 7054 3722 7118 3830
rect 7212 3722 7276 3830
rect 7370 3722 7434 3830
rect 7528 3722 7592 3830
rect 7686 3722 7750 3830
rect 7844 3722 7908 3830
rect 8002 3722 8066 3830
rect 8160 3722 8224 3830
rect 8318 3722 8382 3830
rect 8476 3722 8540 3830
rect 8634 3722 8698 3830
rect 8792 3722 8856 3830
rect 8950 3722 9014 3830
rect 9108 3722 9172 3830
rect 9266 3722 9330 3830
rect 9424 3722 9488 3830
rect 9582 3722 9646 3830
rect 9740 3722 9804 3830
rect 9898 3722 9962 3830
rect 10056 3722 10120 3830
rect 10214 3722 10278 3830
rect 10372 3722 10436 3830
rect 10530 3722 10594 3830
rect 10688 3722 10752 3830
rect 10846 3722 10910 3830
rect 11004 3722 11068 3830
rect 11162 3722 11226 3830
rect 11320 3722 11384 3830
rect 11478 3722 11542 3830
rect 11636 3722 11700 3830
rect 11794 3722 11858 3830
rect 11952 3722 12016 3830
rect 12110 3722 12174 3830
rect 12268 3722 12332 3830
rect 12426 3722 12490 3830
rect 12584 3722 12648 3830
rect 12742 3722 12806 3830
rect 98 3712 172 3722
rect 98 2934 108 3712
rect 164 2934 172 3712
rect 98 2924 172 2934
rect 256 3712 328 3722
rect 256 2930 266 3712
rect 322 2930 328 3712
rect 102 2812 166 2924
rect 256 2920 328 2930
rect 412 3712 488 3722
rect 412 2930 422 3712
rect 478 2930 488 3712
rect 412 2920 488 2930
rect 572 3712 644 3722
rect 572 2930 582 3712
rect 638 2930 644 3712
rect 572 2920 644 2930
rect 728 3712 804 3722
rect 728 2930 738 3712
rect 794 2930 804 3712
rect 728 2920 804 2930
rect 888 3712 960 3722
rect 888 2930 898 3712
rect 954 2930 960 3712
rect 888 2920 960 2930
rect 1044 3712 1120 3722
rect 1044 2930 1054 3712
rect 1110 2930 1120 3712
rect 1044 2920 1120 2930
rect 1204 3712 1276 3722
rect 1204 2930 1214 3712
rect 1270 2930 1276 3712
rect 1204 2920 1276 2930
rect 1360 3712 1436 3722
rect 1360 2930 1370 3712
rect 1426 2930 1436 3712
rect 1360 2920 1436 2930
rect 1520 3712 1592 3722
rect 1520 2930 1530 3712
rect 1586 2930 1592 3712
rect 1520 2920 1592 2930
rect 1676 3712 1752 3722
rect 1676 2930 1686 3712
rect 1742 2930 1752 3712
rect 1676 2920 1752 2930
rect 1836 3712 1908 3722
rect 1836 2930 1846 3712
rect 1902 2930 1908 3712
rect 1836 2920 1908 2930
rect 1992 3712 2068 3722
rect 1992 2930 2002 3712
rect 2058 2930 2068 3712
rect 1992 2920 2068 2930
rect 2152 3712 2224 3722
rect 2152 2930 2162 3712
rect 2218 2930 2224 3712
rect 2152 2920 2224 2930
rect 2308 3712 2384 3722
rect 2308 2930 2318 3712
rect 2374 2930 2384 3712
rect 2308 2920 2384 2930
rect 2468 3712 2540 3722
rect 2468 2930 2478 3712
rect 2534 2930 2540 3712
rect 2468 2920 2540 2930
rect 2624 3712 2700 3722
rect 2624 2930 2634 3712
rect 2690 2930 2700 3712
rect 2624 2920 2700 2930
rect 2784 3712 2856 3722
rect 2784 2930 2794 3712
rect 2850 2930 2856 3712
rect 2784 2920 2856 2930
rect 2940 3712 3016 3722
rect 2940 2930 2950 3712
rect 3006 2930 3016 3712
rect 2940 2920 3016 2930
rect 3100 3712 3172 3722
rect 3100 2930 3110 3712
rect 3166 2930 3172 3712
rect 3100 2920 3172 2930
rect 3256 3712 3332 3722
rect 3256 2930 3266 3712
rect 3322 2930 3332 3712
rect 3256 2920 3332 2930
rect 3416 3712 3488 3722
rect 3416 2930 3426 3712
rect 3482 2930 3488 3712
rect 3416 2920 3488 2930
rect 3572 3712 3648 3722
rect 3572 2930 3582 3712
rect 3638 2930 3648 3712
rect 3572 2920 3648 2930
rect 3732 3712 3804 3722
rect 3732 2930 3742 3712
rect 3798 2930 3804 3712
rect 3732 2920 3804 2930
rect 3888 3712 3964 3722
rect 3888 2930 3898 3712
rect 3954 2930 3964 3712
rect 3888 2920 3964 2930
rect 4048 3712 4120 3722
rect 4048 2930 4058 3712
rect 4114 2930 4120 3712
rect 4048 2920 4120 2930
rect 4204 3712 4280 3722
rect 4204 2930 4214 3712
rect 4270 2930 4280 3712
rect 4204 2920 4280 2930
rect 4364 3712 4436 3722
rect 4364 2930 4374 3712
rect 4430 2930 4436 3712
rect 4364 2920 4436 2930
rect 4520 3712 4596 3722
rect 4520 2930 4530 3712
rect 4586 2930 4596 3712
rect 4520 2920 4596 2930
rect 4680 3712 4752 3722
rect 4680 2930 4690 3712
rect 4746 2930 4752 3712
rect 4680 2920 4752 2930
rect 4836 3712 4912 3722
rect 4836 2930 4846 3712
rect 4902 2930 4912 3712
rect 4836 2920 4912 2930
rect 4996 3712 5068 3722
rect 4996 2930 5006 3712
rect 5062 2930 5068 3712
rect 4996 2920 5068 2930
rect 5152 3712 5228 3722
rect 5152 2930 5162 3712
rect 5218 2930 5228 3712
rect 5152 2920 5228 2930
rect 5312 3712 5384 3722
rect 5312 2930 5322 3712
rect 5378 2930 5384 3712
rect 5312 2920 5384 2930
rect 5468 3712 5544 3722
rect 5468 2930 5478 3712
rect 5534 2930 5544 3712
rect 5468 2920 5544 2930
rect 5628 3712 5700 3722
rect 5628 2930 5638 3712
rect 5694 2930 5700 3712
rect 5628 2920 5700 2930
rect 5784 3712 5860 3722
rect 5784 2930 5794 3712
rect 5850 2930 5860 3712
rect 5784 2920 5860 2930
rect 5944 3712 6016 3722
rect 5944 2930 5954 3712
rect 6010 2930 6016 3712
rect 5944 2920 6016 2930
rect 6100 3712 6176 3722
rect 6100 2930 6110 3712
rect 6166 2930 6176 3712
rect 6100 2920 6176 2930
rect 6260 3712 6332 3722
rect 6260 2930 6270 3712
rect 6326 2930 6332 3712
rect 6260 2920 6332 2930
rect 6416 3712 6492 3722
rect 6416 2930 6426 3712
rect 6482 2930 6492 3712
rect 6416 2920 6492 2930
rect 6576 3712 6648 3722
rect 6576 2930 6586 3712
rect 6642 2930 6648 3712
rect 6576 2920 6648 2930
rect 6732 3712 6808 3722
rect 6732 2930 6742 3712
rect 6798 2930 6808 3712
rect 6732 2920 6808 2930
rect 6892 3712 6964 3722
rect 6892 2930 6902 3712
rect 6958 2930 6964 3712
rect 6892 2920 6964 2930
rect 7048 3712 7124 3722
rect 7048 2930 7058 3712
rect 7114 2930 7124 3712
rect 7048 2920 7124 2930
rect 7208 3712 7280 3722
rect 7208 2930 7218 3712
rect 7274 2930 7280 3712
rect 7208 2920 7280 2930
rect 7364 3712 7440 3722
rect 7364 2930 7374 3712
rect 7430 2930 7440 3712
rect 7364 2920 7440 2930
rect 7524 3712 7596 3722
rect 7524 2930 7534 3712
rect 7590 2930 7596 3712
rect 7524 2920 7596 2930
rect 7680 3712 7756 3722
rect 7680 2930 7690 3712
rect 7746 2930 7756 3712
rect 7680 2920 7756 2930
rect 7840 3712 7912 3722
rect 7840 2930 7850 3712
rect 7906 2930 7912 3712
rect 7840 2920 7912 2930
rect 7996 3712 8072 3722
rect 7996 2930 8006 3712
rect 8062 2930 8072 3712
rect 7996 2920 8072 2930
rect 8156 3712 8228 3722
rect 8156 2930 8166 3712
rect 8222 2930 8228 3712
rect 8156 2920 8228 2930
rect 8312 3712 8388 3722
rect 8312 2930 8322 3712
rect 8378 2930 8388 3712
rect 8312 2920 8388 2930
rect 8472 3712 8544 3722
rect 8472 2930 8482 3712
rect 8538 2930 8544 3712
rect 8472 2920 8544 2930
rect 8628 3712 8704 3722
rect 8628 2930 8638 3712
rect 8694 2930 8704 3712
rect 8628 2920 8704 2930
rect 8788 3712 8860 3722
rect 8788 2930 8798 3712
rect 8854 2930 8860 3712
rect 8788 2920 8860 2930
rect 8944 3712 9020 3722
rect 8944 2930 8954 3712
rect 9010 2930 9020 3712
rect 8944 2920 9020 2930
rect 9104 3712 9176 3722
rect 9104 2930 9114 3712
rect 9170 2930 9176 3712
rect 9104 2920 9176 2930
rect 9260 3712 9336 3722
rect 9260 2930 9270 3712
rect 9326 2930 9336 3712
rect 9260 2920 9336 2930
rect 9420 3712 9492 3722
rect 9420 2930 9430 3712
rect 9486 2930 9492 3712
rect 9420 2920 9492 2930
rect 9576 3712 9652 3722
rect 9576 2930 9586 3712
rect 9642 2930 9652 3712
rect 9576 2920 9652 2930
rect 9736 3712 9808 3722
rect 9736 2930 9746 3712
rect 9802 2930 9808 3712
rect 9736 2920 9808 2930
rect 9892 3712 9968 3722
rect 9892 2930 9902 3712
rect 9958 2930 9968 3712
rect 9892 2920 9968 2930
rect 10052 3712 10124 3722
rect 10052 2930 10062 3712
rect 10118 2930 10124 3712
rect 10052 2920 10124 2930
rect 10208 3712 10284 3722
rect 10208 2930 10218 3712
rect 10274 2930 10284 3712
rect 10208 2920 10284 2930
rect 10368 3712 10440 3722
rect 10368 2930 10378 3712
rect 10434 2930 10440 3712
rect 10368 2920 10440 2930
rect 10524 3712 10600 3722
rect 10524 2930 10534 3712
rect 10590 2930 10600 3712
rect 10524 2920 10600 2930
rect 10684 3712 10756 3722
rect 10684 2930 10694 3712
rect 10750 2930 10756 3712
rect 10684 2920 10756 2930
rect 10840 3712 10916 3722
rect 10840 2930 10850 3712
rect 10906 2930 10916 3712
rect 10840 2920 10916 2930
rect 11000 3712 11072 3722
rect 11000 2930 11010 3712
rect 11066 2930 11072 3712
rect 11000 2920 11072 2930
rect 11156 3712 11232 3722
rect 11156 2930 11166 3712
rect 11222 2930 11232 3712
rect 11156 2920 11232 2930
rect 11316 3712 11388 3722
rect 11316 2930 11326 3712
rect 11382 2930 11388 3712
rect 11316 2920 11388 2930
rect 11472 3712 11548 3722
rect 11472 2930 11482 3712
rect 11538 2930 11548 3712
rect 11472 2920 11548 2930
rect 11632 3712 11704 3722
rect 11632 2930 11642 3712
rect 11698 2930 11704 3712
rect 11632 2920 11704 2930
rect 11788 3712 11864 3722
rect 11788 2930 11798 3712
rect 11854 2930 11864 3712
rect 11788 2920 11864 2930
rect 11948 3712 12020 3722
rect 11948 2930 11958 3712
rect 12014 2930 12020 3712
rect 11948 2920 12020 2930
rect 12104 3712 12180 3722
rect 12104 2930 12114 3712
rect 12170 2930 12180 3712
rect 12104 2920 12180 2930
rect 12264 3712 12336 3722
rect 12264 2930 12274 3712
rect 12330 2930 12336 3712
rect 12264 2920 12336 2930
rect 12420 3712 12496 3722
rect 12420 2930 12430 3712
rect 12486 2930 12496 3712
rect 12420 2920 12496 2930
rect 12580 3712 12652 3722
rect 12580 2930 12590 3712
rect 12646 2930 12652 3712
rect 12580 2920 12652 2930
rect 12736 3712 12812 3722
rect 12736 2930 12746 3712
rect 12802 2930 12812 3712
rect 12736 2920 12812 2930
rect 260 2812 324 2920
rect 418 2812 482 2920
rect 576 2812 640 2920
rect 734 2812 798 2920
rect 892 2812 956 2920
rect 1050 2812 1114 2920
rect 1208 2812 1272 2920
rect 1366 2812 1430 2920
rect 1524 2812 1588 2920
rect 1682 2812 1746 2920
rect 1840 2812 1904 2920
rect 1998 2812 2062 2920
rect 2156 2812 2220 2920
rect 2314 2812 2378 2920
rect 2472 2812 2536 2920
rect 2630 2812 2694 2920
rect 2788 2812 2852 2920
rect 2946 2812 3010 2920
rect 3104 2812 3168 2920
rect 3262 2812 3326 2920
rect 3420 2812 3484 2920
rect 3578 2812 3642 2920
rect 3736 2812 3800 2920
rect 3894 2812 3958 2920
rect 4052 2812 4116 2920
rect 4210 2812 4274 2920
rect 4368 2812 4432 2920
rect 4526 2812 4590 2920
rect 4684 2812 4748 2920
rect 4842 2812 4906 2920
rect 5000 2812 5064 2920
rect 5158 2812 5222 2920
rect 5316 2812 5380 2920
rect 5474 2812 5538 2920
rect 5632 2812 5696 2920
rect 5790 2812 5854 2920
rect 5948 2812 6012 2920
rect 6106 2812 6170 2920
rect 6264 2812 6328 2920
rect 6422 2812 6486 2920
rect 6580 2812 6644 2920
rect 6738 2812 6802 2920
rect 6896 2812 6960 2920
rect 7054 2812 7118 2920
rect 7212 2812 7276 2920
rect 7370 2812 7434 2920
rect 7528 2812 7592 2920
rect 7686 2812 7750 2920
rect 7844 2812 7908 2920
rect 8002 2812 8066 2920
rect 8160 2812 8224 2920
rect 8318 2812 8382 2920
rect 8476 2812 8540 2920
rect 8634 2812 8698 2920
rect 8792 2812 8856 2920
rect 8950 2812 9014 2920
rect 9108 2812 9172 2920
rect 9266 2812 9330 2920
rect 9424 2812 9488 2920
rect 9582 2812 9646 2920
rect 9740 2812 9804 2920
rect 9898 2812 9962 2920
rect 10056 2812 10120 2920
rect 10214 2812 10278 2920
rect 10372 2812 10436 2920
rect 10530 2812 10594 2920
rect 10688 2812 10752 2920
rect 10846 2812 10910 2920
rect 11004 2812 11068 2920
rect 11162 2812 11226 2920
rect 11320 2812 11384 2920
rect 11478 2812 11542 2920
rect 11636 2812 11700 2920
rect 11794 2812 11858 2920
rect 11952 2812 12016 2920
rect 12110 2812 12174 2920
rect 12268 2812 12332 2920
rect 12426 2812 12490 2920
rect 12584 2812 12648 2920
rect 12742 2812 12806 2920
rect 98 2802 172 2812
rect 98 2024 108 2802
rect 164 2024 172 2802
rect 98 2014 172 2024
rect 256 2802 328 2812
rect 256 2020 266 2802
rect 322 2020 328 2802
rect 102 1902 166 2014
rect 256 2010 328 2020
rect 412 2802 488 2812
rect 412 2020 422 2802
rect 478 2020 488 2802
rect 412 2010 488 2020
rect 572 2802 644 2812
rect 572 2020 582 2802
rect 638 2020 644 2802
rect 572 2010 644 2020
rect 728 2802 804 2812
rect 728 2020 738 2802
rect 794 2020 804 2802
rect 728 2010 804 2020
rect 888 2802 960 2812
rect 888 2020 898 2802
rect 954 2020 960 2802
rect 888 2010 960 2020
rect 1044 2802 1120 2812
rect 1044 2020 1054 2802
rect 1110 2020 1120 2802
rect 1044 2010 1120 2020
rect 1204 2802 1276 2812
rect 1204 2020 1214 2802
rect 1270 2020 1276 2802
rect 1204 2010 1276 2020
rect 1360 2802 1436 2812
rect 1360 2020 1370 2802
rect 1426 2020 1436 2802
rect 1360 2010 1436 2020
rect 1520 2802 1592 2812
rect 1520 2020 1530 2802
rect 1586 2020 1592 2802
rect 1520 2010 1592 2020
rect 1676 2802 1752 2812
rect 1676 2020 1686 2802
rect 1742 2020 1752 2802
rect 1676 2010 1752 2020
rect 1836 2802 1908 2812
rect 1836 2020 1846 2802
rect 1902 2020 1908 2802
rect 1836 2010 1908 2020
rect 1992 2802 2068 2812
rect 1992 2020 2002 2802
rect 2058 2020 2068 2802
rect 1992 2010 2068 2020
rect 2152 2802 2224 2812
rect 2152 2020 2162 2802
rect 2218 2020 2224 2802
rect 2152 2010 2224 2020
rect 2308 2802 2384 2812
rect 2308 2020 2318 2802
rect 2374 2020 2384 2802
rect 2308 2010 2384 2020
rect 2468 2802 2540 2812
rect 2468 2020 2478 2802
rect 2534 2020 2540 2802
rect 2468 2010 2540 2020
rect 2624 2802 2700 2812
rect 2624 2020 2634 2802
rect 2690 2020 2700 2802
rect 2624 2010 2700 2020
rect 2784 2802 2856 2812
rect 2784 2020 2794 2802
rect 2850 2020 2856 2802
rect 2784 2010 2856 2020
rect 2940 2802 3016 2812
rect 2940 2020 2950 2802
rect 3006 2020 3016 2802
rect 2940 2010 3016 2020
rect 3100 2802 3172 2812
rect 3100 2020 3110 2802
rect 3166 2020 3172 2802
rect 3100 2010 3172 2020
rect 3256 2802 3332 2812
rect 3256 2020 3266 2802
rect 3322 2020 3332 2802
rect 3256 2010 3332 2020
rect 3416 2802 3488 2812
rect 3416 2020 3426 2802
rect 3482 2020 3488 2802
rect 3416 2010 3488 2020
rect 3572 2802 3648 2812
rect 3572 2020 3582 2802
rect 3638 2020 3648 2802
rect 3572 2010 3648 2020
rect 3732 2802 3804 2812
rect 3732 2020 3742 2802
rect 3798 2020 3804 2802
rect 3732 2010 3804 2020
rect 3888 2802 3964 2812
rect 3888 2020 3898 2802
rect 3954 2020 3964 2802
rect 3888 2010 3964 2020
rect 4048 2802 4120 2812
rect 4048 2020 4058 2802
rect 4114 2020 4120 2802
rect 4048 2010 4120 2020
rect 4204 2802 4280 2812
rect 4204 2020 4214 2802
rect 4270 2020 4280 2802
rect 4204 2010 4280 2020
rect 4364 2802 4436 2812
rect 4364 2020 4374 2802
rect 4430 2020 4436 2802
rect 4364 2010 4436 2020
rect 4520 2802 4596 2812
rect 4520 2020 4530 2802
rect 4586 2020 4596 2802
rect 4520 2010 4596 2020
rect 4680 2802 4752 2812
rect 4680 2020 4690 2802
rect 4746 2020 4752 2802
rect 4680 2010 4752 2020
rect 4836 2802 4912 2812
rect 4836 2020 4846 2802
rect 4902 2020 4912 2802
rect 4836 2010 4912 2020
rect 4996 2802 5068 2812
rect 4996 2020 5006 2802
rect 5062 2020 5068 2802
rect 4996 2010 5068 2020
rect 5152 2802 5228 2812
rect 5152 2020 5162 2802
rect 5218 2020 5228 2802
rect 5152 2010 5228 2020
rect 5312 2802 5384 2812
rect 5312 2020 5322 2802
rect 5378 2020 5384 2802
rect 5312 2010 5384 2020
rect 5468 2802 5544 2812
rect 5468 2020 5478 2802
rect 5534 2020 5544 2802
rect 5468 2010 5544 2020
rect 5628 2802 5700 2812
rect 5628 2020 5638 2802
rect 5694 2020 5700 2802
rect 5628 2010 5700 2020
rect 5784 2802 5860 2812
rect 5784 2020 5794 2802
rect 5850 2020 5860 2802
rect 5784 2010 5860 2020
rect 5944 2802 6016 2812
rect 5944 2020 5954 2802
rect 6010 2020 6016 2802
rect 5944 2010 6016 2020
rect 6100 2802 6176 2812
rect 6100 2020 6110 2802
rect 6166 2020 6176 2802
rect 6100 2010 6176 2020
rect 6260 2802 6332 2812
rect 6260 2020 6270 2802
rect 6326 2020 6332 2802
rect 6260 2010 6332 2020
rect 6416 2802 6492 2812
rect 6416 2020 6426 2802
rect 6482 2020 6492 2802
rect 6416 2010 6492 2020
rect 6576 2802 6648 2812
rect 6576 2020 6586 2802
rect 6642 2020 6648 2802
rect 6576 2010 6648 2020
rect 6732 2802 6808 2812
rect 6732 2020 6742 2802
rect 6798 2020 6808 2802
rect 6732 2010 6808 2020
rect 6892 2802 6964 2812
rect 6892 2020 6902 2802
rect 6958 2020 6964 2802
rect 6892 2010 6964 2020
rect 7048 2802 7124 2812
rect 7048 2020 7058 2802
rect 7114 2020 7124 2802
rect 7048 2010 7124 2020
rect 7208 2802 7280 2812
rect 7208 2020 7218 2802
rect 7274 2020 7280 2802
rect 7208 2010 7280 2020
rect 7364 2802 7440 2812
rect 7364 2020 7374 2802
rect 7430 2020 7440 2802
rect 7364 2010 7440 2020
rect 7524 2802 7596 2812
rect 7524 2020 7534 2802
rect 7590 2020 7596 2802
rect 7524 2010 7596 2020
rect 7680 2802 7756 2812
rect 7680 2020 7690 2802
rect 7746 2020 7756 2802
rect 7680 2010 7756 2020
rect 7840 2802 7912 2812
rect 7840 2020 7850 2802
rect 7906 2020 7912 2802
rect 7840 2010 7912 2020
rect 7996 2802 8072 2812
rect 7996 2020 8006 2802
rect 8062 2020 8072 2802
rect 7996 2010 8072 2020
rect 8156 2802 8228 2812
rect 8156 2020 8166 2802
rect 8222 2020 8228 2802
rect 8156 2010 8228 2020
rect 8312 2802 8388 2812
rect 8312 2020 8322 2802
rect 8378 2020 8388 2802
rect 8312 2010 8388 2020
rect 8472 2802 8544 2812
rect 8472 2020 8482 2802
rect 8538 2020 8544 2802
rect 8472 2010 8544 2020
rect 8628 2802 8704 2812
rect 8628 2020 8638 2802
rect 8694 2020 8704 2802
rect 8628 2010 8704 2020
rect 8788 2802 8860 2812
rect 8788 2020 8798 2802
rect 8854 2020 8860 2802
rect 8788 2010 8860 2020
rect 8944 2802 9020 2812
rect 8944 2020 8954 2802
rect 9010 2020 9020 2802
rect 8944 2010 9020 2020
rect 9104 2802 9176 2812
rect 9104 2020 9114 2802
rect 9170 2020 9176 2802
rect 9104 2010 9176 2020
rect 9260 2802 9336 2812
rect 9260 2020 9270 2802
rect 9326 2020 9336 2802
rect 9260 2010 9336 2020
rect 9420 2802 9492 2812
rect 9420 2020 9430 2802
rect 9486 2020 9492 2802
rect 9420 2010 9492 2020
rect 9576 2802 9652 2812
rect 9576 2020 9586 2802
rect 9642 2020 9652 2802
rect 9576 2010 9652 2020
rect 9736 2802 9808 2812
rect 9736 2020 9746 2802
rect 9802 2020 9808 2802
rect 9736 2010 9808 2020
rect 9892 2802 9968 2812
rect 9892 2020 9902 2802
rect 9958 2020 9968 2802
rect 9892 2010 9968 2020
rect 10052 2802 10124 2812
rect 10052 2020 10062 2802
rect 10118 2020 10124 2802
rect 10052 2010 10124 2020
rect 10208 2802 10284 2812
rect 10208 2020 10218 2802
rect 10274 2020 10284 2802
rect 10208 2010 10284 2020
rect 10368 2802 10440 2812
rect 10368 2020 10378 2802
rect 10434 2020 10440 2802
rect 10368 2010 10440 2020
rect 10524 2802 10600 2812
rect 10524 2020 10534 2802
rect 10590 2020 10600 2802
rect 10524 2010 10600 2020
rect 10684 2802 10756 2812
rect 10684 2020 10694 2802
rect 10750 2020 10756 2802
rect 10684 2010 10756 2020
rect 10840 2802 10916 2812
rect 10840 2020 10850 2802
rect 10906 2020 10916 2802
rect 10840 2010 10916 2020
rect 11000 2802 11072 2812
rect 11000 2020 11010 2802
rect 11066 2020 11072 2802
rect 11000 2010 11072 2020
rect 11156 2802 11232 2812
rect 11156 2020 11166 2802
rect 11222 2020 11232 2802
rect 11156 2010 11232 2020
rect 11316 2802 11388 2812
rect 11316 2020 11326 2802
rect 11382 2020 11388 2802
rect 11316 2010 11388 2020
rect 11472 2802 11548 2812
rect 11472 2020 11482 2802
rect 11538 2020 11548 2802
rect 11472 2010 11548 2020
rect 11632 2802 11704 2812
rect 11632 2020 11642 2802
rect 11698 2020 11704 2802
rect 11632 2010 11704 2020
rect 11788 2802 11864 2812
rect 11788 2020 11798 2802
rect 11854 2020 11864 2802
rect 11788 2010 11864 2020
rect 11948 2802 12020 2812
rect 11948 2020 11958 2802
rect 12014 2020 12020 2802
rect 11948 2010 12020 2020
rect 12104 2802 12180 2812
rect 12104 2020 12114 2802
rect 12170 2020 12180 2802
rect 12104 2010 12180 2020
rect 12264 2802 12336 2812
rect 12264 2020 12274 2802
rect 12330 2020 12336 2802
rect 12264 2010 12336 2020
rect 12420 2802 12496 2812
rect 12420 2020 12430 2802
rect 12486 2020 12496 2802
rect 12420 2010 12496 2020
rect 12580 2802 12652 2812
rect 12580 2020 12590 2802
rect 12646 2020 12652 2802
rect 12580 2010 12652 2020
rect 12736 2802 12812 2812
rect 12736 2020 12746 2802
rect 12802 2020 12812 2802
rect 12736 2010 12812 2020
rect 260 1902 324 2010
rect 418 1902 482 2010
rect 576 1902 640 2010
rect 734 1902 798 2010
rect 892 1902 956 2010
rect 1050 1902 1114 2010
rect 1208 1902 1272 2010
rect 1366 1902 1430 2010
rect 1524 1902 1588 2010
rect 1682 1902 1746 2010
rect 1840 1902 1904 2010
rect 1998 1902 2062 2010
rect 2156 1902 2220 2010
rect 2314 1902 2378 2010
rect 2472 1902 2536 2010
rect 2630 1902 2694 2010
rect 2788 1902 2852 2010
rect 2946 1902 3010 2010
rect 3104 1902 3168 2010
rect 3262 1902 3326 2010
rect 3420 1902 3484 2010
rect 3578 1902 3642 2010
rect 3736 1902 3800 2010
rect 3894 1902 3958 2010
rect 4052 1902 4116 2010
rect 4210 1902 4274 2010
rect 4368 1902 4432 2010
rect 4526 1902 4590 2010
rect 4684 1902 4748 2010
rect 4842 1902 4906 2010
rect 5000 1902 5064 2010
rect 5158 1902 5222 2010
rect 5316 1902 5380 2010
rect 5474 1902 5538 2010
rect 5632 1902 5696 2010
rect 5790 1902 5854 2010
rect 5948 1902 6012 2010
rect 6106 1902 6170 2010
rect 6264 1902 6328 2010
rect 6422 1902 6486 2010
rect 6580 1902 6644 2010
rect 6738 1902 6802 2010
rect 6896 1902 6960 2010
rect 7054 1902 7118 2010
rect 7212 1902 7276 2010
rect 7370 1902 7434 2010
rect 7528 1902 7592 2010
rect 7686 1902 7750 2010
rect 7844 1902 7908 2010
rect 8002 1902 8066 2010
rect 8160 1902 8224 2010
rect 8318 1902 8382 2010
rect 8476 1902 8540 2010
rect 8634 1902 8698 2010
rect 8792 1902 8856 2010
rect 8950 1902 9014 2010
rect 9108 1902 9172 2010
rect 9266 1902 9330 2010
rect 9424 1902 9488 2010
rect 9582 1902 9646 2010
rect 9740 1902 9804 2010
rect 9898 1902 9962 2010
rect 10056 1902 10120 2010
rect 10214 1902 10278 2010
rect 10372 1902 10436 2010
rect 10530 1902 10594 2010
rect 10688 1902 10752 2010
rect 10846 1902 10910 2010
rect 11004 1902 11068 2010
rect 11162 1902 11226 2010
rect 11320 1902 11384 2010
rect 11478 1902 11542 2010
rect 11636 1902 11700 2010
rect 11794 1902 11858 2010
rect 11952 1902 12016 2010
rect 12110 1902 12174 2010
rect 12268 1902 12332 2010
rect 12426 1902 12490 2010
rect 12584 1902 12648 2010
rect 12742 1902 12806 2010
rect 98 1892 172 1902
rect 98 1114 108 1892
rect 164 1114 172 1892
rect 98 1104 172 1114
rect 256 1892 328 1902
rect 256 1110 266 1892
rect 322 1110 328 1892
rect 102 992 166 1104
rect 256 1100 328 1110
rect 412 1892 488 1902
rect 412 1110 422 1892
rect 478 1110 488 1892
rect 412 1100 488 1110
rect 572 1892 644 1902
rect 572 1110 582 1892
rect 638 1110 644 1892
rect 572 1100 644 1110
rect 728 1892 804 1902
rect 728 1110 738 1892
rect 794 1110 804 1892
rect 728 1100 804 1110
rect 888 1892 960 1902
rect 888 1110 898 1892
rect 954 1110 960 1892
rect 888 1100 960 1110
rect 1044 1892 1120 1902
rect 1044 1110 1054 1892
rect 1110 1110 1120 1892
rect 1044 1100 1120 1110
rect 1204 1892 1276 1902
rect 1204 1110 1214 1892
rect 1270 1110 1276 1892
rect 1204 1100 1276 1110
rect 1360 1892 1436 1902
rect 1360 1110 1370 1892
rect 1426 1110 1436 1892
rect 1360 1100 1436 1110
rect 1520 1892 1592 1902
rect 1520 1110 1530 1892
rect 1586 1110 1592 1892
rect 1520 1100 1592 1110
rect 1676 1892 1752 1902
rect 1676 1110 1686 1892
rect 1742 1110 1752 1892
rect 1676 1100 1752 1110
rect 1836 1892 1908 1902
rect 1836 1110 1846 1892
rect 1902 1110 1908 1892
rect 1836 1100 1908 1110
rect 1992 1892 2068 1902
rect 1992 1110 2002 1892
rect 2058 1110 2068 1892
rect 1992 1100 2068 1110
rect 2152 1892 2224 1902
rect 2152 1110 2162 1892
rect 2218 1110 2224 1892
rect 2152 1100 2224 1110
rect 2308 1892 2384 1902
rect 2308 1110 2318 1892
rect 2374 1110 2384 1892
rect 2308 1100 2384 1110
rect 2468 1892 2540 1902
rect 2468 1110 2478 1892
rect 2534 1110 2540 1892
rect 2468 1100 2540 1110
rect 2624 1892 2700 1902
rect 2624 1110 2634 1892
rect 2690 1110 2700 1892
rect 2624 1100 2700 1110
rect 2784 1892 2856 1902
rect 2784 1110 2794 1892
rect 2850 1110 2856 1892
rect 2784 1100 2856 1110
rect 2940 1892 3016 1902
rect 2940 1110 2950 1892
rect 3006 1110 3016 1892
rect 2940 1100 3016 1110
rect 3100 1892 3172 1902
rect 3100 1110 3110 1892
rect 3166 1110 3172 1892
rect 3100 1100 3172 1110
rect 3256 1892 3332 1902
rect 3256 1110 3266 1892
rect 3322 1110 3332 1892
rect 3256 1100 3332 1110
rect 3416 1892 3488 1902
rect 3416 1110 3426 1892
rect 3482 1110 3488 1892
rect 3416 1100 3488 1110
rect 3572 1892 3648 1902
rect 3572 1110 3582 1892
rect 3638 1110 3648 1892
rect 3572 1100 3648 1110
rect 3732 1892 3804 1902
rect 3732 1110 3742 1892
rect 3798 1110 3804 1892
rect 3732 1100 3804 1110
rect 3888 1892 3964 1902
rect 3888 1110 3898 1892
rect 3954 1110 3964 1892
rect 3888 1100 3964 1110
rect 4048 1892 4120 1902
rect 4048 1110 4058 1892
rect 4114 1110 4120 1892
rect 4048 1100 4120 1110
rect 4204 1892 4280 1902
rect 4204 1110 4214 1892
rect 4270 1110 4280 1892
rect 4204 1100 4280 1110
rect 4364 1892 4436 1902
rect 4364 1110 4374 1892
rect 4430 1110 4436 1892
rect 4364 1100 4436 1110
rect 4520 1892 4596 1902
rect 4520 1110 4530 1892
rect 4586 1110 4596 1892
rect 4520 1100 4596 1110
rect 4680 1892 4752 1902
rect 4680 1110 4690 1892
rect 4746 1110 4752 1892
rect 4680 1100 4752 1110
rect 4836 1892 4912 1902
rect 4836 1110 4846 1892
rect 4902 1110 4912 1892
rect 4836 1100 4912 1110
rect 4996 1892 5068 1902
rect 4996 1110 5006 1892
rect 5062 1110 5068 1892
rect 4996 1100 5068 1110
rect 5152 1892 5228 1902
rect 5152 1110 5162 1892
rect 5218 1110 5228 1892
rect 5152 1100 5228 1110
rect 5312 1892 5384 1902
rect 5312 1110 5322 1892
rect 5378 1110 5384 1892
rect 5312 1100 5384 1110
rect 5468 1892 5544 1902
rect 5468 1110 5478 1892
rect 5534 1110 5544 1892
rect 5468 1100 5544 1110
rect 5628 1892 5700 1902
rect 5628 1110 5638 1892
rect 5694 1110 5700 1892
rect 5628 1100 5700 1110
rect 5784 1892 5860 1902
rect 5784 1110 5794 1892
rect 5850 1110 5860 1892
rect 5784 1100 5860 1110
rect 5944 1892 6016 1902
rect 5944 1110 5954 1892
rect 6010 1110 6016 1892
rect 5944 1100 6016 1110
rect 6100 1892 6176 1902
rect 6100 1110 6110 1892
rect 6166 1110 6176 1892
rect 6100 1100 6176 1110
rect 6260 1892 6332 1902
rect 6260 1110 6270 1892
rect 6326 1110 6332 1892
rect 6260 1100 6332 1110
rect 6416 1892 6492 1902
rect 6416 1110 6426 1892
rect 6482 1110 6492 1892
rect 6416 1100 6492 1110
rect 6576 1892 6648 1902
rect 6576 1110 6586 1892
rect 6642 1110 6648 1892
rect 6576 1100 6648 1110
rect 6732 1892 6808 1902
rect 6732 1110 6742 1892
rect 6798 1110 6808 1892
rect 6732 1100 6808 1110
rect 6892 1892 6964 1902
rect 6892 1110 6902 1892
rect 6958 1110 6964 1892
rect 6892 1100 6964 1110
rect 7048 1892 7124 1902
rect 7048 1110 7058 1892
rect 7114 1110 7124 1892
rect 7048 1100 7124 1110
rect 7208 1892 7280 1902
rect 7208 1110 7218 1892
rect 7274 1110 7280 1892
rect 7208 1100 7280 1110
rect 7364 1892 7440 1902
rect 7364 1110 7374 1892
rect 7430 1110 7440 1892
rect 7364 1100 7440 1110
rect 7524 1892 7596 1902
rect 7524 1110 7534 1892
rect 7590 1110 7596 1892
rect 7524 1100 7596 1110
rect 7680 1892 7756 1902
rect 7680 1110 7690 1892
rect 7746 1110 7756 1892
rect 7680 1100 7756 1110
rect 7840 1892 7912 1902
rect 7840 1110 7850 1892
rect 7906 1110 7912 1892
rect 7840 1100 7912 1110
rect 7996 1892 8072 1902
rect 7996 1110 8006 1892
rect 8062 1110 8072 1892
rect 7996 1100 8072 1110
rect 8156 1892 8228 1902
rect 8156 1110 8166 1892
rect 8222 1110 8228 1892
rect 8156 1100 8228 1110
rect 8312 1892 8388 1902
rect 8312 1110 8322 1892
rect 8378 1110 8388 1892
rect 8312 1100 8388 1110
rect 8472 1892 8544 1902
rect 8472 1110 8482 1892
rect 8538 1110 8544 1892
rect 8472 1100 8544 1110
rect 8628 1892 8704 1902
rect 8628 1110 8638 1892
rect 8694 1110 8704 1892
rect 8628 1100 8704 1110
rect 8788 1892 8860 1902
rect 8788 1110 8798 1892
rect 8854 1110 8860 1892
rect 8788 1100 8860 1110
rect 8944 1892 9020 1902
rect 8944 1110 8954 1892
rect 9010 1110 9020 1892
rect 8944 1100 9020 1110
rect 9104 1892 9176 1902
rect 9104 1110 9114 1892
rect 9170 1110 9176 1892
rect 9104 1100 9176 1110
rect 9260 1892 9336 1902
rect 9260 1110 9270 1892
rect 9326 1110 9336 1892
rect 9260 1100 9336 1110
rect 9420 1892 9492 1902
rect 9420 1110 9430 1892
rect 9486 1110 9492 1892
rect 9420 1100 9492 1110
rect 9576 1892 9652 1902
rect 9576 1110 9586 1892
rect 9642 1110 9652 1892
rect 9576 1100 9652 1110
rect 9736 1892 9808 1902
rect 9736 1110 9746 1892
rect 9802 1110 9808 1892
rect 9736 1100 9808 1110
rect 9892 1892 9968 1902
rect 9892 1110 9902 1892
rect 9958 1110 9968 1892
rect 9892 1100 9968 1110
rect 10052 1892 10124 1902
rect 10052 1110 10062 1892
rect 10118 1110 10124 1892
rect 10052 1100 10124 1110
rect 10208 1892 10284 1902
rect 10208 1110 10218 1892
rect 10274 1110 10284 1892
rect 10208 1100 10284 1110
rect 10368 1892 10440 1902
rect 10368 1110 10378 1892
rect 10434 1110 10440 1892
rect 10368 1100 10440 1110
rect 10524 1892 10600 1902
rect 10524 1110 10534 1892
rect 10590 1110 10600 1892
rect 10524 1100 10600 1110
rect 10684 1892 10756 1902
rect 10684 1110 10694 1892
rect 10750 1110 10756 1892
rect 10684 1100 10756 1110
rect 10840 1892 10916 1902
rect 10840 1110 10850 1892
rect 10906 1110 10916 1892
rect 10840 1100 10916 1110
rect 11000 1892 11072 1902
rect 11000 1110 11010 1892
rect 11066 1110 11072 1892
rect 11000 1100 11072 1110
rect 11156 1892 11232 1902
rect 11156 1110 11166 1892
rect 11222 1110 11232 1892
rect 11156 1100 11232 1110
rect 11316 1892 11388 1902
rect 11316 1110 11326 1892
rect 11382 1110 11388 1892
rect 11316 1100 11388 1110
rect 11472 1892 11548 1902
rect 11472 1110 11482 1892
rect 11538 1110 11548 1892
rect 11472 1100 11548 1110
rect 11632 1892 11704 1902
rect 11632 1110 11642 1892
rect 11698 1110 11704 1892
rect 11632 1100 11704 1110
rect 11788 1892 11864 1902
rect 11788 1110 11798 1892
rect 11854 1110 11864 1892
rect 11788 1100 11864 1110
rect 11948 1892 12020 1902
rect 11948 1110 11958 1892
rect 12014 1110 12020 1892
rect 11948 1100 12020 1110
rect 12104 1892 12180 1902
rect 12104 1110 12114 1892
rect 12170 1110 12180 1892
rect 12104 1100 12180 1110
rect 12264 1892 12336 1902
rect 12264 1110 12274 1892
rect 12330 1110 12336 1892
rect 12264 1100 12336 1110
rect 12420 1892 12496 1902
rect 12420 1110 12430 1892
rect 12486 1110 12496 1892
rect 12420 1100 12496 1110
rect 12580 1892 12652 1902
rect 12580 1110 12590 1892
rect 12646 1110 12652 1892
rect 12580 1100 12652 1110
rect 12736 1892 12812 1902
rect 12736 1110 12746 1892
rect 12802 1110 12812 1892
rect 12736 1100 12812 1110
rect 260 992 324 1100
rect 418 992 482 1100
rect 576 992 640 1100
rect 734 992 798 1100
rect 892 992 956 1100
rect 1050 992 1114 1100
rect 1208 992 1272 1100
rect 1366 992 1430 1100
rect 1524 992 1588 1100
rect 1682 992 1746 1100
rect 1840 992 1904 1100
rect 1998 992 2062 1100
rect 2156 992 2220 1100
rect 2314 992 2378 1100
rect 2472 992 2536 1100
rect 2630 992 2694 1100
rect 2788 992 2852 1100
rect 2946 992 3010 1100
rect 3104 992 3168 1100
rect 3262 992 3326 1100
rect 3420 992 3484 1100
rect 3578 992 3642 1100
rect 3736 992 3800 1100
rect 3894 992 3958 1100
rect 4052 992 4116 1100
rect 4210 992 4274 1100
rect 4368 992 4432 1100
rect 4526 992 4590 1100
rect 4684 992 4748 1100
rect 4842 992 4906 1100
rect 5000 992 5064 1100
rect 5158 992 5222 1100
rect 5316 992 5380 1100
rect 5474 992 5538 1100
rect 5632 992 5696 1100
rect 5790 992 5854 1100
rect 5948 992 6012 1100
rect 6106 992 6170 1100
rect 6264 992 6328 1100
rect 6422 992 6486 1100
rect 6580 992 6644 1100
rect 6738 992 6802 1100
rect 6896 992 6960 1100
rect 7054 992 7118 1100
rect 7212 992 7276 1100
rect 7370 992 7434 1100
rect 7528 992 7592 1100
rect 7686 992 7750 1100
rect 7844 992 7908 1100
rect 8002 992 8066 1100
rect 8160 992 8224 1100
rect 8318 992 8382 1100
rect 8476 992 8540 1100
rect 8634 992 8698 1100
rect 8792 992 8856 1100
rect 8950 992 9014 1100
rect 9108 992 9172 1100
rect 9266 992 9330 1100
rect 9424 992 9488 1100
rect 9582 992 9646 1100
rect 9740 992 9804 1100
rect 9898 992 9962 1100
rect 10056 992 10120 1100
rect 10214 992 10278 1100
rect 10372 992 10436 1100
rect 10530 992 10594 1100
rect 10688 992 10752 1100
rect 10846 992 10910 1100
rect 11004 992 11068 1100
rect 11162 992 11226 1100
rect 11320 992 11384 1100
rect 11478 992 11542 1100
rect 11636 992 11700 1100
rect 11794 992 11858 1100
rect 11952 992 12016 1100
rect 12110 992 12174 1100
rect 12268 992 12332 1100
rect 12426 992 12490 1100
rect 12584 992 12648 1100
rect 12742 992 12806 1100
rect 98 982 172 992
rect 98 204 108 982
rect 164 204 172 982
rect 98 194 172 204
rect 256 982 328 992
rect 256 200 266 982
rect 322 200 328 982
rect 102 -66 166 194
rect 256 190 328 200
rect 412 982 488 992
rect 412 200 422 982
rect 478 200 488 982
rect 412 190 488 200
rect 572 982 644 992
rect 572 200 582 982
rect 638 200 644 982
rect 572 190 644 200
rect 728 982 804 992
rect 728 200 738 982
rect 794 200 804 982
rect 728 190 804 200
rect 888 982 960 992
rect 888 200 898 982
rect 954 200 960 982
rect 888 190 960 200
rect 1044 982 1120 992
rect 1044 200 1054 982
rect 1110 200 1120 982
rect 1044 190 1120 200
rect 1204 982 1276 992
rect 1204 200 1214 982
rect 1270 200 1276 982
rect 1204 190 1276 200
rect 1360 982 1436 992
rect 1360 200 1370 982
rect 1426 200 1436 982
rect 1360 190 1436 200
rect 1520 982 1592 992
rect 1520 200 1530 982
rect 1586 200 1592 982
rect 1520 190 1592 200
rect 1676 982 1752 992
rect 1676 200 1686 982
rect 1742 200 1752 982
rect 1676 190 1752 200
rect 1836 982 1908 992
rect 1836 200 1846 982
rect 1902 200 1908 982
rect 1836 190 1908 200
rect 1992 982 2068 992
rect 1992 200 2002 982
rect 2058 200 2068 982
rect 1992 190 2068 200
rect 2152 982 2224 992
rect 2152 200 2162 982
rect 2218 200 2224 982
rect 2152 190 2224 200
rect 2308 982 2384 992
rect 2308 200 2318 982
rect 2374 200 2384 982
rect 2308 190 2384 200
rect 2468 982 2540 992
rect 2468 200 2478 982
rect 2534 200 2540 982
rect 2468 190 2540 200
rect 2624 982 2700 992
rect 2624 200 2634 982
rect 2690 200 2700 982
rect 2624 190 2700 200
rect 2784 982 2856 992
rect 2784 200 2794 982
rect 2850 200 2856 982
rect 2784 190 2856 200
rect 2940 982 3016 992
rect 2940 200 2950 982
rect 3006 200 3016 982
rect 2940 190 3016 200
rect 3100 982 3172 992
rect 3100 200 3110 982
rect 3166 200 3172 982
rect 3100 190 3172 200
rect 3256 982 3332 992
rect 3256 200 3266 982
rect 3322 200 3332 982
rect 3256 190 3332 200
rect 3416 982 3488 992
rect 3416 200 3426 982
rect 3482 200 3488 982
rect 3416 190 3488 200
rect 3572 982 3648 992
rect 3572 200 3582 982
rect 3638 200 3648 982
rect 3572 190 3648 200
rect 3732 982 3804 992
rect 3732 200 3742 982
rect 3798 200 3804 982
rect 3732 190 3804 200
rect 3888 982 3964 992
rect 3888 200 3898 982
rect 3954 200 3964 982
rect 3888 190 3964 200
rect 4048 982 4120 992
rect 4048 200 4058 982
rect 4114 200 4120 982
rect 4048 190 4120 200
rect 4204 982 4280 992
rect 4204 200 4214 982
rect 4270 200 4280 982
rect 4204 190 4280 200
rect 4364 982 4436 992
rect 4364 200 4374 982
rect 4430 200 4436 982
rect 4364 190 4436 200
rect 4520 982 4596 992
rect 4520 200 4530 982
rect 4586 200 4596 982
rect 4520 190 4596 200
rect 4680 982 4752 992
rect 4680 200 4690 982
rect 4746 200 4752 982
rect 4680 190 4752 200
rect 4836 982 4912 992
rect 4836 200 4846 982
rect 4902 200 4912 982
rect 4836 190 4912 200
rect 4996 982 5068 992
rect 4996 200 5006 982
rect 5062 200 5068 982
rect 4996 190 5068 200
rect 5152 982 5228 992
rect 5152 200 5162 982
rect 5218 200 5228 982
rect 5152 190 5228 200
rect 5312 982 5384 992
rect 5312 200 5322 982
rect 5378 200 5384 982
rect 5312 190 5384 200
rect 5468 982 5544 992
rect 5468 200 5478 982
rect 5534 200 5544 982
rect 5468 190 5544 200
rect 5628 982 5700 992
rect 5628 200 5638 982
rect 5694 200 5700 982
rect 5628 190 5700 200
rect 5784 982 5860 992
rect 5784 200 5794 982
rect 5850 200 5860 982
rect 5784 190 5860 200
rect 5944 982 6016 992
rect 5944 200 5954 982
rect 6010 200 6016 982
rect 5944 190 6016 200
rect 6100 982 6176 992
rect 6100 200 6110 982
rect 6166 200 6176 982
rect 6100 190 6176 200
rect 6260 982 6332 992
rect 6260 200 6270 982
rect 6326 200 6332 982
rect 6260 190 6332 200
rect 6416 982 6492 992
rect 6416 200 6426 982
rect 6482 200 6492 982
rect 6416 190 6492 200
rect 6576 982 6648 992
rect 6576 200 6586 982
rect 6642 200 6648 982
rect 6576 190 6648 200
rect 6732 982 6808 992
rect 6732 200 6742 982
rect 6798 200 6808 982
rect 6732 190 6808 200
rect 6892 982 6964 992
rect 6892 200 6902 982
rect 6958 200 6964 982
rect 6892 190 6964 200
rect 7048 982 7124 992
rect 7048 200 7058 982
rect 7114 200 7124 982
rect 7048 190 7124 200
rect 7208 982 7280 992
rect 7208 200 7218 982
rect 7274 200 7280 982
rect 7208 190 7280 200
rect 7364 982 7440 992
rect 7364 200 7374 982
rect 7430 200 7440 982
rect 7364 190 7440 200
rect 7524 982 7596 992
rect 7524 200 7534 982
rect 7590 200 7596 982
rect 7524 190 7596 200
rect 7680 982 7756 992
rect 7680 200 7690 982
rect 7746 200 7756 982
rect 7680 190 7756 200
rect 7840 982 7912 992
rect 7840 200 7850 982
rect 7906 200 7912 982
rect 7840 190 7912 200
rect 7996 982 8072 992
rect 7996 200 8006 982
rect 8062 200 8072 982
rect 7996 190 8072 200
rect 8156 982 8228 992
rect 8156 200 8166 982
rect 8222 200 8228 982
rect 8156 190 8228 200
rect 8312 982 8388 992
rect 8312 200 8322 982
rect 8378 200 8388 982
rect 8312 190 8388 200
rect 8472 982 8544 992
rect 8472 200 8482 982
rect 8538 200 8544 982
rect 8472 190 8544 200
rect 8628 982 8704 992
rect 8628 200 8638 982
rect 8694 200 8704 982
rect 8628 190 8704 200
rect 8788 982 8860 992
rect 8788 200 8798 982
rect 8854 200 8860 982
rect 8788 190 8860 200
rect 8944 982 9020 992
rect 8944 200 8954 982
rect 9010 200 9020 982
rect 8944 190 9020 200
rect 9104 982 9176 992
rect 9104 200 9114 982
rect 9170 200 9176 982
rect 9104 190 9176 200
rect 9260 982 9336 992
rect 9260 200 9270 982
rect 9326 200 9336 982
rect 9260 190 9336 200
rect 9420 982 9492 992
rect 9420 200 9430 982
rect 9486 200 9492 982
rect 9420 190 9492 200
rect 9576 982 9652 992
rect 9576 200 9586 982
rect 9642 200 9652 982
rect 9576 190 9652 200
rect 9736 982 9808 992
rect 9736 200 9746 982
rect 9802 200 9808 982
rect 9736 190 9808 200
rect 9892 982 9968 992
rect 9892 200 9902 982
rect 9958 200 9968 982
rect 9892 190 9968 200
rect 10052 982 10124 992
rect 10052 200 10062 982
rect 10118 200 10124 982
rect 10052 190 10124 200
rect 10208 982 10284 992
rect 10208 200 10218 982
rect 10274 200 10284 982
rect 10208 190 10284 200
rect 10368 982 10440 992
rect 10368 200 10378 982
rect 10434 200 10440 982
rect 10368 190 10440 200
rect 10524 982 10600 992
rect 10524 200 10534 982
rect 10590 200 10600 982
rect 10524 190 10600 200
rect 10684 982 10756 992
rect 10684 200 10694 982
rect 10750 200 10756 982
rect 10684 190 10756 200
rect 10840 982 10916 992
rect 10840 200 10850 982
rect 10906 200 10916 982
rect 10840 190 10916 200
rect 11000 982 11072 992
rect 11000 200 11010 982
rect 11066 200 11072 982
rect 11000 190 11072 200
rect 11156 982 11232 992
rect 11156 200 11166 982
rect 11222 200 11232 982
rect 11156 190 11232 200
rect 11316 982 11388 992
rect 11316 200 11326 982
rect 11382 200 11388 982
rect 11316 190 11388 200
rect 11472 982 11548 992
rect 11472 200 11482 982
rect 11538 200 11548 982
rect 11472 190 11548 200
rect 11632 982 11704 992
rect 11632 200 11642 982
rect 11698 200 11704 982
rect 11632 190 11704 200
rect 11788 982 11864 992
rect 11788 200 11798 982
rect 11854 200 11864 982
rect 11788 190 11864 200
rect 11948 982 12020 992
rect 11948 200 11958 982
rect 12014 200 12020 982
rect 11948 190 12020 200
rect 12104 982 12180 992
rect 12104 200 12114 982
rect 12170 200 12180 982
rect 12104 190 12180 200
rect 12264 982 12336 992
rect 12264 200 12274 982
rect 12330 200 12336 982
rect 12264 190 12336 200
rect 12420 982 12496 992
rect 12420 200 12430 982
rect 12486 200 12496 982
rect 12420 190 12496 200
rect 12580 982 12652 992
rect 12580 200 12590 982
rect 12646 200 12652 982
rect 12580 190 12652 200
rect 12736 982 12812 992
rect 12736 200 12746 982
rect 12802 200 12812 982
rect 12736 190 12812 200
rect 260 -66 324 190
rect 418 -66 482 190
rect 576 -66 640 190
rect 734 -66 798 190
rect 892 -66 956 190
rect 1050 -66 1114 190
rect 1208 -66 1272 190
rect 1366 -66 1430 190
rect 1524 -66 1588 190
rect 1682 -66 1746 190
rect 1840 -66 1904 190
rect 1998 -66 2062 190
rect 2156 -66 2220 190
rect 2314 -66 2378 190
rect 2472 -66 2536 190
rect 2630 -66 2694 190
rect 2788 -66 2852 190
rect 2946 -66 3010 190
rect 3104 -66 3168 190
rect 3262 -66 3326 190
rect 3420 -66 3484 190
rect 3578 -66 3642 190
rect 3736 -66 3800 190
rect 3894 -66 3958 190
rect 4052 -66 4116 190
rect 4210 -66 4274 190
rect 4368 -66 4432 190
rect 4526 -66 4590 190
rect 4684 -66 4748 190
rect 4842 -66 4906 190
rect 5000 -66 5064 190
rect 5158 -66 5222 190
rect 5316 -66 5380 190
rect 5474 -66 5538 190
rect 5632 -66 5696 190
rect 5790 -66 5854 190
rect 5948 -66 6012 190
rect 6106 -66 6170 190
rect 6264 -66 6328 190
rect 6422 -66 6486 190
rect 6580 -66 6644 190
rect 6738 -66 6802 190
rect 6896 -66 6960 190
rect 7054 -66 7118 190
rect 7212 -66 7276 190
rect 7370 -66 7434 190
rect 7528 -66 7592 190
rect 7686 -66 7750 190
rect 7844 -66 7908 190
rect 8002 -66 8066 190
rect 8160 -66 8224 190
rect 8318 -66 8382 190
rect 8476 -66 8540 190
rect 8634 -66 8698 190
rect 8792 -66 8856 190
rect 8950 -66 9014 190
rect 9108 -66 9172 190
rect 9266 -66 9330 190
rect 9424 -66 9488 190
rect 9582 -66 9646 190
rect 9740 -66 9804 190
rect 9898 -66 9962 190
rect 10056 -66 10120 190
rect 10214 -66 10278 190
rect 10372 -66 10436 190
rect 10530 -66 10594 190
rect 10688 -66 10752 190
rect 10846 -66 10910 190
rect 11004 -66 11068 190
rect 11162 -66 11226 190
rect 11320 -66 11384 190
rect 11478 -66 11542 190
rect 11636 -66 11700 190
rect 11794 -66 11858 190
rect 11952 -66 12016 190
rect 12110 -66 12174 190
rect 12268 -66 12332 190
rect 12426 -66 12490 190
rect 12584 -66 12648 190
rect 12742 -66 12806 190
use sky130_fd_pr__nfet_g5v0d10v5_KBPKF4  sky130_fd_pr__nfet_g5v0d10v5_KBPKF4_0
timestamp 1664842101
transform 1 0 6453 0 1 2412
box -6519 -2478 6519 2478
<< end >>
