magic
tech sky130A
timestamp 1667507583
<< nwell >>
rect -10470 -698 10470 698
<< pwell >>
rect -10560 698 10560 788
rect -10560 -698 -10470 698
rect 10470 -698 10560 698
rect -10560 -788 10560 -698
<< mvpsubdiff >>
rect -10542 764 10542 770
rect -10542 747 -10488 764
rect 10488 747 10542 764
rect -10542 741 10542 747
rect -10542 716 -10513 741
rect -10542 -716 -10536 716
rect -10519 -716 -10513 716
rect 10513 716 10542 741
rect -10542 -741 -10513 -716
rect 10513 -716 10519 716
rect 10536 -716 10542 716
rect 10513 -741 10542 -716
rect -10542 -747 10542 -741
rect -10542 -764 -10488 -747
rect 10488 -764 10542 -747
rect -10542 -770 10542 -764
<< mvnsubdiff >>
rect -10437 659 -9805 665
rect -10437 642 -10383 659
rect -9859 642 -9805 659
rect -10437 636 -9805 642
rect -10437 611 -10408 636
rect -10437 87 -10431 611
rect -10414 87 -10408 611
rect -9834 611 -9805 636
rect -10437 62 -10408 87
rect -9834 87 -9828 611
rect -9811 87 -9805 611
rect -9834 62 -9805 87
rect -10437 56 -9805 62
rect -10437 39 -10383 56
rect -9859 39 -9805 56
rect -10437 33 -9805 39
rect -9739 659 -9107 665
rect -9739 642 -9685 659
rect -9161 642 -9107 659
rect -9739 636 -9107 642
rect -9739 611 -9710 636
rect -9739 87 -9733 611
rect -9716 87 -9710 611
rect -9136 611 -9107 636
rect -9739 62 -9710 87
rect -9136 87 -9130 611
rect -9113 87 -9107 611
rect -9136 62 -9107 87
rect -9739 56 -9107 62
rect -9739 39 -9685 56
rect -9161 39 -9107 56
rect -9739 33 -9107 39
rect -9041 659 -8409 665
rect -9041 642 -8987 659
rect -8463 642 -8409 659
rect -9041 636 -8409 642
rect -9041 611 -9012 636
rect -9041 87 -9035 611
rect -9018 87 -9012 611
rect -8438 611 -8409 636
rect -9041 62 -9012 87
rect -8438 87 -8432 611
rect -8415 87 -8409 611
rect -8438 62 -8409 87
rect -9041 56 -8409 62
rect -9041 39 -8987 56
rect -8463 39 -8409 56
rect -9041 33 -8409 39
rect -8343 659 -7711 665
rect -8343 642 -8289 659
rect -7765 642 -7711 659
rect -8343 636 -7711 642
rect -8343 611 -8314 636
rect -8343 87 -8337 611
rect -8320 87 -8314 611
rect -7740 611 -7711 636
rect -8343 62 -8314 87
rect -7740 87 -7734 611
rect -7717 87 -7711 611
rect -7740 62 -7711 87
rect -8343 56 -7711 62
rect -8343 39 -8289 56
rect -7765 39 -7711 56
rect -8343 33 -7711 39
rect -7645 659 -7013 665
rect -7645 642 -7591 659
rect -7067 642 -7013 659
rect -7645 636 -7013 642
rect -7645 611 -7616 636
rect -7645 87 -7639 611
rect -7622 87 -7616 611
rect -7042 611 -7013 636
rect -7645 62 -7616 87
rect -7042 87 -7036 611
rect -7019 87 -7013 611
rect -7042 62 -7013 87
rect -7645 56 -7013 62
rect -7645 39 -7591 56
rect -7067 39 -7013 56
rect -7645 33 -7013 39
rect -6947 659 -6315 665
rect -6947 642 -6893 659
rect -6369 642 -6315 659
rect -6947 636 -6315 642
rect -6947 611 -6918 636
rect -6947 87 -6941 611
rect -6924 87 -6918 611
rect -6344 611 -6315 636
rect -6947 62 -6918 87
rect -6344 87 -6338 611
rect -6321 87 -6315 611
rect -6344 62 -6315 87
rect -6947 56 -6315 62
rect -6947 39 -6893 56
rect -6369 39 -6315 56
rect -6947 33 -6315 39
rect -6249 659 -5617 665
rect -6249 642 -6195 659
rect -5671 642 -5617 659
rect -6249 636 -5617 642
rect -6249 611 -6220 636
rect -6249 87 -6243 611
rect -6226 87 -6220 611
rect -5646 611 -5617 636
rect -6249 62 -6220 87
rect -5646 87 -5640 611
rect -5623 87 -5617 611
rect -5646 62 -5617 87
rect -6249 56 -5617 62
rect -6249 39 -6195 56
rect -5671 39 -5617 56
rect -6249 33 -5617 39
rect -5551 659 -4919 665
rect -5551 642 -5497 659
rect -4973 642 -4919 659
rect -5551 636 -4919 642
rect -5551 611 -5522 636
rect -5551 87 -5545 611
rect -5528 87 -5522 611
rect -4948 611 -4919 636
rect -5551 62 -5522 87
rect -4948 87 -4942 611
rect -4925 87 -4919 611
rect -4948 62 -4919 87
rect -5551 56 -4919 62
rect -5551 39 -5497 56
rect -4973 39 -4919 56
rect -5551 33 -4919 39
rect -4853 659 -4221 665
rect -4853 642 -4799 659
rect -4275 642 -4221 659
rect -4853 636 -4221 642
rect -4853 611 -4824 636
rect -4853 87 -4847 611
rect -4830 87 -4824 611
rect -4250 611 -4221 636
rect -4853 62 -4824 87
rect -4250 87 -4244 611
rect -4227 87 -4221 611
rect -4250 62 -4221 87
rect -4853 56 -4221 62
rect -4853 39 -4799 56
rect -4275 39 -4221 56
rect -4853 33 -4221 39
rect -4155 659 -3523 665
rect -4155 642 -4101 659
rect -3577 642 -3523 659
rect -4155 636 -3523 642
rect -4155 611 -4126 636
rect -4155 87 -4149 611
rect -4132 87 -4126 611
rect -3552 611 -3523 636
rect -4155 62 -4126 87
rect -3552 87 -3546 611
rect -3529 87 -3523 611
rect -3552 62 -3523 87
rect -4155 56 -3523 62
rect -4155 39 -4101 56
rect -3577 39 -3523 56
rect -4155 33 -3523 39
rect -3457 659 -2825 665
rect -3457 642 -3403 659
rect -2879 642 -2825 659
rect -3457 636 -2825 642
rect -3457 611 -3428 636
rect -3457 87 -3451 611
rect -3434 87 -3428 611
rect -2854 611 -2825 636
rect -3457 62 -3428 87
rect -2854 87 -2848 611
rect -2831 87 -2825 611
rect -2854 62 -2825 87
rect -3457 56 -2825 62
rect -3457 39 -3403 56
rect -2879 39 -2825 56
rect -3457 33 -2825 39
rect -2759 659 -2127 665
rect -2759 642 -2705 659
rect -2181 642 -2127 659
rect -2759 636 -2127 642
rect -2759 611 -2730 636
rect -2759 87 -2753 611
rect -2736 87 -2730 611
rect -2156 611 -2127 636
rect -2759 62 -2730 87
rect -2156 87 -2150 611
rect -2133 87 -2127 611
rect -2156 62 -2127 87
rect -2759 56 -2127 62
rect -2759 39 -2705 56
rect -2181 39 -2127 56
rect -2759 33 -2127 39
rect -2061 659 -1429 665
rect -2061 642 -2007 659
rect -1483 642 -1429 659
rect -2061 636 -1429 642
rect -2061 611 -2032 636
rect -2061 87 -2055 611
rect -2038 87 -2032 611
rect -1458 611 -1429 636
rect -2061 62 -2032 87
rect -1458 87 -1452 611
rect -1435 87 -1429 611
rect -1458 62 -1429 87
rect -2061 56 -1429 62
rect -2061 39 -2007 56
rect -1483 39 -1429 56
rect -2061 33 -1429 39
rect -1363 659 -731 665
rect -1363 642 -1309 659
rect -785 642 -731 659
rect -1363 636 -731 642
rect -1363 611 -1334 636
rect -1363 87 -1357 611
rect -1340 87 -1334 611
rect -760 611 -731 636
rect -1363 62 -1334 87
rect -760 87 -754 611
rect -737 87 -731 611
rect -760 62 -731 87
rect -1363 56 -731 62
rect -1363 39 -1309 56
rect -785 39 -731 56
rect -1363 33 -731 39
rect -665 659 -33 665
rect -665 642 -611 659
rect -87 642 -33 659
rect -665 636 -33 642
rect -665 611 -636 636
rect -665 87 -659 611
rect -642 87 -636 611
rect -62 611 -33 636
rect -665 62 -636 87
rect -62 87 -56 611
rect -39 87 -33 611
rect -62 62 -33 87
rect -665 56 -33 62
rect -665 39 -611 56
rect -87 39 -33 56
rect -665 33 -33 39
rect 33 659 665 665
rect 33 642 87 659
rect 611 642 665 659
rect 33 636 665 642
rect 33 611 62 636
rect 33 87 39 611
rect 56 87 62 611
rect 636 611 665 636
rect 33 62 62 87
rect 636 87 642 611
rect 659 87 665 611
rect 636 62 665 87
rect 33 56 665 62
rect 33 39 87 56
rect 611 39 665 56
rect 33 33 665 39
rect 731 659 1363 665
rect 731 642 785 659
rect 1309 642 1363 659
rect 731 636 1363 642
rect 731 611 760 636
rect 731 87 737 611
rect 754 87 760 611
rect 1334 611 1363 636
rect 731 62 760 87
rect 1334 87 1340 611
rect 1357 87 1363 611
rect 1334 62 1363 87
rect 731 56 1363 62
rect 731 39 785 56
rect 1309 39 1363 56
rect 731 33 1363 39
rect 1429 659 2061 665
rect 1429 642 1483 659
rect 2007 642 2061 659
rect 1429 636 2061 642
rect 1429 611 1458 636
rect 1429 87 1435 611
rect 1452 87 1458 611
rect 2032 611 2061 636
rect 1429 62 1458 87
rect 2032 87 2038 611
rect 2055 87 2061 611
rect 2032 62 2061 87
rect 1429 56 2061 62
rect 1429 39 1483 56
rect 2007 39 2061 56
rect 1429 33 2061 39
rect 2127 659 2759 665
rect 2127 642 2181 659
rect 2705 642 2759 659
rect 2127 636 2759 642
rect 2127 611 2156 636
rect 2127 87 2133 611
rect 2150 87 2156 611
rect 2730 611 2759 636
rect 2127 62 2156 87
rect 2730 87 2736 611
rect 2753 87 2759 611
rect 2730 62 2759 87
rect 2127 56 2759 62
rect 2127 39 2181 56
rect 2705 39 2759 56
rect 2127 33 2759 39
rect 2825 659 3457 665
rect 2825 642 2879 659
rect 3403 642 3457 659
rect 2825 636 3457 642
rect 2825 611 2854 636
rect 2825 87 2831 611
rect 2848 87 2854 611
rect 3428 611 3457 636
rect 2825 62 2854 87
rect 3428 87 3434 611
rect 3451 87 3457 611
rect 3428 62 3457 87
rect 2825 56 3457 62
rect 2825 39 2879 56
rect 3403 39 3457 56
rect 2825 33 3457 39
rect 3523 659 4155 665
rect 3523 642 3577 659
rect 4101 642 4155 659
rect 3523 636 4155 642
rect 3523 611 3552 636
rect 3523 87 3529 611
rect 3546 87 3552 611
rect 4126 611 4155 636
rect 3523 62 3552 87
rect 4126 87 4132 611
rect 4149 87 4155 611
rect 4126 62 4155 87
rect 3523 56 4155 62
rect 3523 39 3577 56
rect 4101 39 4155 56
rect 3523 33 4155 39
rect 4221 659 4853 665
rect 4221 642 4275 659
rect 4799 642 4853 659
rect 4221 636 4853 642
rect 4221 611 4250 636
rect 4221 87 4227 611
rect 4244 87 4250 611
rect 4824 611 4853 636
rect 4221 62 4250 87
rect 4824 87 4830 611
rect 4847 87 4853 611
rect 4824 62 4853 87
rect 4221 56 4853 62
rect 4221 39 4275 56
rect 4799 39 4853 56
rect 4221 33 4853 39
rect 4919 659 5551 665
rect 4919 642 4973 659
rect 5497 642 5551 659
rect 4919 636 5551 642
rect 4919 611 4948 636
rect 4919 87 4925 611
rect 4942 87 4948 611
rect 5522 611 5551 636
rect 4919 62 4948 87
rect 5522 87 5528 611
rect 5545 87 5551 611
rect 5522 62 5551 87
rect 4919 56 5551 62
rect 4919 39 4973 56
rect 5497 39 5551 56
rect 4919 33 5551 39
rect 5617 659 6249 665
rect 5617 642 5671 659
rect 6195 642 6249 659
rect 5617 636 6249 642
rect 5617 611 5646 636
rect 5617 87 5623 611
rect 5640 87 5646 611
rect 6220 611 6249 636
rect 5617 62 5646 87
rect 6220 87 6226 611
rect 6243 87 6249 611
rect 6220 62 6249 87
rect 5617 56 6249 62
rect 5617 39 5671 56
rect 6195 39 6249 56
rect 5617 33 6249 39
rect 6315 659 6947 665
rect 6315 642 6369 659
rect 6893 642 6947 659
rect 6315 636 6947 642
rect 6315 611 6344 636
rect 6315 87 6321 611
rect 6338 87 6344 611
rect 6918 611 6947 636
rect 6315 62 6344 87
rect 6918 87 6924 611
rect 6941 87 6947 611
rect 6918 62 6947 87
rect 6315 56 6947 62
rect 6315 39 6369 56
rect 6893 39 6947 56
rect 6315 33 6947 39
rect 7013 659 7645 665
rect 7013 642 7067 659
rect 7591 642 7645 659
rect 7013 636 7645 642
rect 7013 611 7042 636
rect 7013 87 7019 611
rect 7036 87 7042 611
rect 7616 611 7645 636
rect 7013 62 7042 87
rect 7616 87 7622 611
rect 7639 87 7645 611
rect 7616 62 7645 87
rect 7013 56 7645 62
rect 7013 39 7067 56
rect 7591 39 7645 56
rect 7013 33 7645 39
rect 7711 659 8343 665
rect 7711 642 7765 659
rect 8289 642 8343 659
rect 7711 636 8343 642
rect 7711 611 7740 636
rect 7711 87 7717 611
rect 7734 87 7740 611
rect 8314 611 8343 636
rect 7711 62 7740 87
rect 8314 87 8320 611
rect 8337 87 8343 611
rect 8314 62 8343 87
rect 7711 56 8343 62
rect 7711 39 7765 56
rect 8289 39 8343 56
rect 7711 33 8343 39
rect 8409 659 9041 665
rect 8409 642 8463 659
rect 8987 642 9041 659
rect 8409 636 9041 642
rect 8409 611 8438 636
rect 8409 87 8415 611
rect 8432 87 8438 611
rect 9012 611 9041 636
rect 8409 62 8438 87
rect 9012 87 9018 611
rect 9035 87 9041 611
rect 9012 62 9041 87
rect 8409 56 9041 62
rect 8409 39 8463 56
rect 8987 39 9041 56
rect 8409 33 9041 39
rect 9107 659 9739 665
rect 9107 642 9161 659
rect 9685 642 9739 659
rect 9107 636 9739 642
rect 9107 611 9136 636
rect 9107 87 9113 611
rect 9130 87 9136 611
rect 9710 611 9739 636
rect 9107 62 9136 87
rect 9710 87 9716 611
rect 9733 87 9739 611
rect 9710 62 9739 87
rect 9107 56 9739 62
rect 9107 39 9161 56
rect 9685 39 9739 56
rect 9107 33 9739 39
rect 9805 659 10437 665
rect 9805 642 9859 659
rect 10383 642 10437 659
rect 9805 636 10437 642
rect 9805 611 9834 636
rect 9805 87 9811 611
rect 9828 87 9834 611
rect 10408 611 10437 636
rect 9805 62 9834 87
rect 10408 87 10414 611
rect 10431 87 10437 611
rect 10408 62 10437 87
rect 9805 56 10437 62
rect 9805 39 9859 56
rect 10383 39 10437 56
rect 9805 33 10437 39
rect -10437 -39 -9805 -33
rect -10437 -56 -10383 -39
rect -9859 -56 -9805 -39
rect -10437 -62 -9805 -56
rect -10437 -87 -10408 -62
rect -10437 -611 -10431 -87
rect -10414 -611 -10408 -87
rect -9834 -87 -9805 -62
rect -10437 -636 -10408 -611
rect -9834 -611 -9828 -87
rect -9811 -611 -9805 -87
rect -9834 -636 -9805 -611
rect -10437 -642 -9805 -636
rect -10437 -659 -10383 -642
rect -9859 -659 -9805 -642
rect -10437 -665 -9805 -659
rect -9739 -39 -9107 -33
rect -9739 -56 -9685 -39
rect -9161 -56 -9107 -39
rect -9739 -62 -9107 -56
rect -9739 -87 -9710 -62
rect -9739 -611 -9733 -87
rect -9716 -611 -9710 -87
rect -9136 -87 -9107 -62
rect -9739 -636 -9710 -611
rect -9136 -611 -9130 -87
rect -9113 -611 -9107 -87
rect -9136 -636 -9107 -611
rect -9739 -642 -9107 -636
rect -9739 -659 -9685 -642
rect -9161 -659 -9107 -642
rect -9739 -665 -9107 -659
rect -9041 -39 -8409 -33
rect -9041 -56 -8987 -39
rect -8463 -56 -8409 -39
rect -9041 -62 -8409 -56
rect -9041 -87 -9012 -62
rect -9041 -611 -9035 -87
rect -9018 -611 -9012 -87
rect -8438 -87 -8409 -62
rect -9041 -636 -9012 -611
rect -8438 -611 -8432 -87
rect -8415 -611 -8409 -87
rect -8438 -636 -8409 -611
rect -9041 -642 -8409 -636
rect -9041 -659 -8987 -642
rect -8463 -659 -8409 -642
rect -9041 -665 -8409 -659
rect -8343 -39 -7711 -33
rect -8343 -56 -8289 -39
rect -7765 -56 -7711 -39
rect -8343 -62 -7711 -56
rect -8343 -87 -8314 -62
rect -8343 -611 -8337 -87
rect -8320 -611 -8314 -87
rect -7740 -87 -7711 -62
rect -8343 -636 -8314 -611
rect -7740 -611 -7734 -87
rect -7717 -611 -7711 -87
rect -7740 -636 -7711 -611
rect -8343 -642 -7711 -636
rect -8343 -659 -8289 -642
rect -7765 -659 -7711 -642
rect -8343 -665 -7711 -659
rect -7645 -39 -7013 -33
rect -7645 -56 -7591 -39
rect -7067 -56 -7013 -39
rect -7645 -62 -7013 -56
rect -7645 -87 -7616 -62
rect -7645 -611 -7639 -87
rect -7622 -611 -7616 -87
rect -7042 -87 -7013 -62
rect -7645 -636 -7616 -611
rect -7042 -611 -7036 -87
rect -7019 -611 -7013 -87
rect -7042 -636 -7013 -611
rect -7645 -642 -7013 -636
rect -7645 -659 -7591 -642
rect -7067 -659 -7013 -642
rect -7645 -665 -7013 -659
rect -6947 -39 -6315 -33
rect -6947 -56 -6893 -39
rect -6369 -56 -6315 -39
rect -6947 -62 -6315 -56
rect -6947 -87 -6918 -62
rect -6947 -611 -6941 -87
rect -6924 -611 -6918 -87
rect -6344 -87 -6315 -62
rect -6947 -636 -6918 -611
rect -6344 -611 -6338 -87
rect -6321 -611 -6315 -87
rect -6344 -636 -6315 -611
rect -6947 -642 -6315 -636
rect -6947 -659 -6893 -642
rect -6369 -659 -6315 -642
rect -6947 -665 -6315 -659
rect -6249 -39 -5617 -33
rect -6249 -56 -6195 -39
rect -5671 -56 -5617 -39
rect -6249 -62 -5617 -56
rect -6249 -87 -6220 -62
rect -6249 -611 -6243 -87
rect -6226 -611 -6220 -87
rect -5646 -87 -5617 -62
rect -6249 -636 -6220 -611
rect -5646 -611 -5640 -87
rect -5623 -611 -5617 -87
rect -5646 -636 -5617 -611
rect -6249 -642 -5617 -636
rect -6249 -659 -6195 -642
rect -5671 -659 -5617 -642
rect -6249 -665 -5617 -659
rect -5551 -39 -4919 -33
rect -5551 -56 -5497 -39
rect -4973 -56 -4919 -39
rect -5551 -62 -4919 -56
rect -5551 -87 -5522 -62
rect -5551 -611 -5545 -87
rect -5528 -611 -5522 -87
rect -4948 -87 -4919 -62
rect -5551 -636 -5522 -611
rect -4948 -611 -4942 -87
rect -4925 -611 -4919 -87
rect -4948 -636 -4919 -611
rect -5551 -642 -4919 -636
rect -5551 -659 -5497 -642
rect -4973 -659 -4919 -642
rect -5551 -665 -4919 -659
rect -4853 -39 -4221 -33
rect -4853 -56 -4799 -39
rect -4275 -56 -4221 -39
rect -4853 -62 -4221 -56
rect -4853 -87 -4824 -62
rect -4853 -611 -4847 -87
rect -4830 -611 -4824 -87
rect -4250 -87 -4221 -62
rect -4853 -636 -4824 -611
rect -4250 -611 -4244 -87
rect -4227 -611 -4221 -87
rect -4250 -636 -4221 -611
rect -4853 -642 -4221 -636
rect -4853 -659 -4799 -642
rect -4275 -659 -4221 -642
rect -4853 -665 -4221 -659
rect -4155 -39 -3523 -33
rect -4155 -56 -4101 -39
rect -3577 -56 -3523 -39
rect -4155 -62 -3523 -56
rect -4155 -87 -4126 -62
rect -4155 -611 -4149 -87
rect -4132 -611 -4126 -87
rect -3552 -87 -3523 -62
rect -4155 -636 -4126 -611
rect -3552 -611 -3546 -87
rect -3529 -611 -3523 -87
rect -3552 -636 -3523 -611
rect -4155 -642 -3523 -636
rect -4155 -659 -4101 -642
rect -3577 -659 -3523 -642
rect -4155 -665 -3523 -659
rect -3457 -39 -2825 -33
rect -3457 -56 -3403 -39
rect -2879 -56 -2825 -39
rect -3457 -62 -2825 -56
rect -3457 -87 -3428 -62
rect -3457 -611 -3451 -87
rect -3434 -611 -3428 -87
rect -2854 -87 -2825 -62
rect -3457 -636 -3428 -611
rect -2854 -611 -2848 -87
rect -2831 -611 -2825 -87
rect -2854 -636 -2825 -611
rect -3457 -642 -2825 -636
rect -3457 -659 -3403 -642
rect -2879 -659 -2825 -642
rect -3457 -665 -2825 -659
rect -2759 -39 -2127 -33
rect -2759 -56 -2705 -39
rect -2181 -56 -2127 -39
rect -2759 -62 -2127 -56
rect -2759 -87 -2730 -62
rect -2759 -611 -2753 -87
rect -2736 -611 -2730 -87
rect -2156 -87 -2127 -62
rect -2759 -636 -2730 -611
rect -2156 -611 -2150 -87
rect -2133 -611 -2127 -87
rect -2156 -636 -2127 -611
rect -2759 -642 -2127 -636
rect -2759 -659 -2705 -642
rect -2181 -659 -2127 -642
rect -2759 -665 -2127 -659
rect -2061 -39 -1429 -33
rect -2061 -56 -2007 -39
rect -1483 -56 -1429 -39
rect -2061 -62 -1429 -56
rect -2061 -87 -2032 -62
rect -2061 -611 -2055 -87
rect -2038 -611 -2032 -87
rect -1458 -87 -1429 -62
rect -2061 -636 -2032 -611
rect -1458 -611 -1452 -87
rect -1435 -611 -1429 -87
rect -1458 -636 -1429 -611
rect -2061 -642 -1429 -636
rect -2061 -659 -2007 -642
rect -1483 -659 -1429 -642
rect -2061 -665 -1429 -659
rect -1363 -39 -731 -33
rect -1363 -56 -1309 -39
rect -785 -56 -731 -39
rect -1363 -62 -731 -56
rect -1363 -87 -1334 -62
rect -1363 -611 -1357 -87
rect -1340 -611 -1334 -87
rect -760 -87 -731 -62
rect -1363 -636 -1334 -611
rect -760 -611 -754 -87
rect -737 -611 -731 -87
rect -760 -636 -731 -611
rect -1363 -642 -731 -636
rect -1363 -659 -1309 -642
rect -785 -659 -731 -642
rect -1363 -665 -731 -659
rect -665 -39 -33 -33
rect -665 -56 -611 -39
rect -87 -56 -33 -39
rect -665 -62 -33 -56
rect -665 -87 -636 -62
rect -665 -611 -659 -87
rect -642 -611 -636 -87
rect -62 -87 -33 -62
rect -665 -636 -636 -611
rect -62 -611 -56 -87
rect -39 -611 -33 -87
rect -62 -636 -33 -611
rect -665 -642 -33 -636
rect -665 -659 -611 -642
rect -87 -659 -33 -642
rect -665 -665 -33 -659
rect 33 -39 665 -33
rect 33 -56 87 -39
rect 611 -56 665 -39
rect 33 -62 665 -56
rect 33 -87 62 -62
rect 33 -611 39 -87
rect 56 -611 62 -87
rect 636 -87 665 -62
rect 33 -636 62 -611
rect 636 -611 642 -87
rect 659 -611 665 -87
rect 636 -636 665 -611
rect 33 -642 665 -636
rect 33 -659 87 -642
rect 611 -659 665 -642
rect 33 -665 665 -659
rect 731 -39 1363 -33
rect 731 -56 785 -39
rect 1309 -56 1363 -39
rect 731 -62 1363 -56
rect 731 -87 760 -62
rect 731 -611 737 -87
rect 754 -611 760 -87
rect 1334 -87 1363 -62
rect 731 -636 760 -611
rect 1334 -611 1340 -87
rect 1357 -611 1363 -87
rect 1334 -636 1363 -611
rect 731 -642 1363 -636
rect 731 -659 785 -642
rect 1309 -659 1363 -642
rect 731 -665 1363 -659
rect 1429 -39 2061 -33
rect 1429 -56 1483 -39
rect 2007 -56 2061 -39
rect 1429 -62 2061 -56
rect 1429 -87 1458 -62
rect 1429 -611 1435 -87
rect 1452 -611 1458 -87
rect 2032 -87 2061 -62
rect 1429 -636 1458 -611
rect 2032 -611 2038 -87
rect 2055 -611 2061 -87
rect 2032 -636 2061 -611
rect 1429 -642 2061 -636
rect 1429 -659 1483 -642
rect 2007 -659 2061 -642
rect 1429 -665 2061 -659
rect 2127 -39 2759 -33
rect 2127 -56 2181 -39
rect 2705 -56 2759 -39
rect 2127 -62 2759 -56
rect 2127 -87 2156 -62
rect 2127 -611 2133 -87
rect 2150 -611 2156 -87
rect 2730 -87 2759 -62
rect 2127 -636 2156 -611
rect 2730 -611 2736 -87
rect 2753 -611 2759 -87
rect 2730 -636 2759 -611
rect 2127 -642 2759 -636
rect 2127 -659 2181 -642
rect 2705 -659 2759 -642
rect 2127 -665 2759 -659
rect 2825 -39 3457 -33
rect 2825 -56 2879 -39
rect 3403 -56 3457 -39
rect 2825 -62 3457 -56
rect 2825 -87 2854 -62
rect 2825 -611 2831 -87
rect 2848 -611 2854 -87
rect 3428 -87 3457 -62
rect 2825 -636 2854 -611
rect 3428 -611 3434 -87
rect 3451 -611 3457 -87
rect 3428 -636 3457 -611
rect 2825 -642 3457 -636
rect 2825 -659 2879 -642
rect 3403 -659 3457 -642
rect 2825 -665 3457 -659
rect 3523 -39 4155 -33
rect 3523 -56 3577 -39
rect 4101 -56 4155 -39
rect 3523 -62 4155 -56
rect 3523 -87 3552 -62
rect 3523 -611 3529 -87
rect 3546 -611 3552 -87
rect 4126 -87 4155 -62
rect 3523 -636 3552 -611
rect 4126 -611 4132 -87
rect 4149 -611 4155 -87
rect 4126 -636 4155 -611
rect 3523 -642 4155 -636
rect 3523 -659 3577 -642
rect 4101 -659 4155 -642
rect 3523 -665 4155 -659
rect 4221 -39 4853 -33
rect 4221 -56 4275 -39
rect 4799 -56 4853 -39
rect 4221 -62 4853 -56
rect 4221 -87 4250 -62
rect 4221 -611 4227 -87
rect 4244 -611 4250 -87
rect 4824 -87 4853 -62
rect 4221 -636 4250 -611
rect 4824 -611 4830 -87
rect 4847 -611 4853 -87
rect 4824 -636 4853 -611
rect 4221 -642 4853 -636
rect 4221 -659 4275 -642
rect 4799 -659 4853 -642
rect 4221 -665 4853 -659
rect 4919 -39 5551 -33
rect 4919 -56 4973 -39
rect 5497 -56 5551 -39
rect 4919 -62 5551 -56
rect 4919 -87 4948 -62
rect 4919 -611 4925 -87
rect 4942 -611 4948 -87
rect 5522 -87 5551 -62
rect 4919 -636 4948 -611
rect 5522 -611 5528 -87
rect 5545 -611 5551 -87
rect 5522 -636 5551 -611
rect 4919 -642 5551 -636
rect 4919 -659 4973 -642
rect 5497 -659 5551 -642
rect 4919 -665 5551 -659
rect 5617 -39 6249 -33
rect 5617 -56 5671 -39
rect 6195 -56 6249 -39
rect 5617 -62 6249 -56
rect 5617 -87 5646 -62
rect 5617 -611 5623 -87
rect 5640 -611 5646 -87
rect 6220 -87 6249 -62
rect 5617 -636 5646 -611
rect 6220 -611 6226 -87
rect 6243 -611 6249 -87
rect 6220 -636 6249 -611
rect 5617 -642 6249 -636
rect 5617 -659 5671 -642
rect 6195 -659 6249 -642
rect 5617 -665 6249 -659
rect 6315 -39 6947 -33
rect 6315 -56 6369 -39
rect 6893 -56 6947 -39
rect 6315 -62 6947 -56
rect 6315 -87 6344 -62
rect 6315 -611 6321 -87
rect 6338 -611 6344 -87
rect 6918 -87 6947 -62
rect 6315 -636 6344 -611
rect 6918 -611 6924 -87
rect 6941 -611 6947 -87
rect 6918 -636 6947 -611
rect 6315 -642 6947 -636
rect 6315 -659 6369 -642
rect 6893 -659 6947 -642
rect 6315 -665 6947 -659
rect 7013 -39 7645 -33
rect 7013 -56 7067 -39
rect 7591 -56 7645 -39
rect 7013 -62 7645 -56
rect 7013 -87 7042 -62
rect 7013 -611 7019 -87
rect 7036 -611 7042 -87
rect 7616 -87 7645 -62
rect 7013 -636 7042 -611
rect 7616 -611 7622 -87
rect 7639 -611 7645 -87
rect 7616 -636 7645 -611
rect 7013 -642 7645 -636
rect 7013 -659 7067 -642
rect 7591 -659 7645 -642
rect 7013 -665 7645 -659
rect 7711 -39 8343 -33
rect 7711 -56 7765 -39
rect 8289 -56 8343 -39
rect 7711 -62 8343 -56
rect 7711 -87 7740 -62
rect 7711 -611 7717 -87
rect 7734 -611 7740 -87
rect 8314 -87 8343 -62
rect 7711 -636 7740 -611
rect 8314 -611 8320 -87
rect 8337 -611 8343 -87
rect 8314 -636 8343 -611
rect 7711 -642 8343 -636
rect 7711 -659 7765 -642
rect 8289 -659 8343 -642
rect 7711 -665 8343 -659
rect 8409 -39 9041 -33
rect 8409 -56 8463 -39
rect 8987 -56 9041 -39
rect 8409 -62 9041 -56
rect 8409 -87 8438 -62
rect 8409 -611 8415 -87
rect 8432 -611 8438 -87
rect 9012 -87 9041 -62
rect 8409 -636 8438 -611
rect 9012 -611 9018 -87
rect 9035 -611 9041 -87
rect 9012 -636 9041 -611
rect 8409 -642 9041 -636
rect 8409 -659 8463 -642
rect 8987 -659 9041 -642
rect 8409 -665 9041 -659
rect 9107 -39 9739 -33
rect 9107 -56 9161 -39
rect 9685 -56 9739 -39
rect 9107 -62 9739 -56
rect 9107 -87 9136 -62
rect 9107 -611 9113 -87
rect 9130 -611 9136 -87
rect 9710 -87 9739 -62
rect 9107 -636 9136 -611
rect 9710 -611 9716 -87
rect 9733 -611 9739 -87
rect 9710 -636 9739 -611
rect 9107 -642 9739 -636
rect 9107 -659 9161 -642
rect 9685 -659 9739 -642
rect 9107 -665 9739 -659
rect 9805 -39 10437 -33
rect 9805 -56 9859 -39
rect 10383 -56 10437 -39
rect 9805 -62 10437 -56
rect 9805 -87 9834 -62
rect 9805 -611 9811 -87
rect 9828 -611 9834 -87
rect 10408 -87 10437 -62
rect 9805 -636 9834 -611
rect 10408 -611 10414 -87
rect 10431 -611 10437 -87
rect 10408 -636 10437 -611
rect 9805 -642 10437 -636
rect 9805 -659 9859 -642
rect 10383 -659 10437 -642
rect 9805 -665 10437 -659
<< mvpsubdiffcont >>
rect -10488 747 10488 764
rect -10536 -716 -10519 716
rect 10519 -716 10536 716
rect -10488 -764 10488 -747
<< mvnsubdiffcont >>
rect -10383 642 -9859 659
rect -10431 87 -10414 611
rect -9828 87 -9811 611
rect -10383 39 -9859 56
rect -9685 642 -9161 659
rect -9733 87 -9716 611
rect -9130 87 -9113 611
rect -9685 39 -9161 56
rect -8987 642 -8463 659
rect -9035 87 -9018 611
rect -8432 87 -8415 611
rect -8987 39 -8463 56
rect -8289 642 -7765 659
rect -8337 87 -8320 611
rect -7734 87 -7717 611
rect -8289 39 -7765 56
rect -7591 642 -7067 659
rect -7639 87 -7622 611
rect -7036 87 -7019 611
rect -7591 39 -7067 56
rect -6893 642 -6369 659
rect -6941 87 -6924 611
rect -6338 87 -6321 611
rect -6893 39 -6369 56
rect -6195 642 -5671 659
rect -6243 87 -6226 611
rect -5640 87 -5623 611
rect -6195 39 -5671 56
rect -5497 642 -4973 659
rect -5545 87 -5528 611
rect -4942 87 -4925 611
rect -5497 39 -4973 56
rect -4799 642 -4275 659
rect -4847 87 -4830 611
rect -4244 87 -4227 611
rect -4799 39 -4275 56
rect -4101 642 -3577 659
rect -4149 87 -4132 611
rect -3546 87 -3529 611
rect -4101 39 -3577 56
rect -3403 642 -2879 659
rect -3451 87 -3434 611
rect -2848 87 -2831 611
rect -3403 39 -2879 56
rect -2705 642 -2181 659
rect -2753 87 -2736 611
rect -2150 87 -2133 611
rect -2705 39 -2181 56
rect -2007 642 -1483 659
rect -2055 87 -2038 611
rect -1452 87 -1435 611
rect -2007 39 -1483 56
rect -1309 642 -785 659
rect -1357 87 -1340 611
rect -754 87 -737 611
rect -1309 39 -785 56
rect -611 642 -87 659
rect -659 87 -642 611
rect -56 87 -39 611
rect -611 39 -87 56
rect 87 642 611 659
rect 39 87 56 611
rect 642 87 659 611
rect 87 39 611 56
rect 785 642 1309 659
rect 737 87 754 611
rect 1340 87 1357 611
rect 785 39 1309 56
rect 1483 642 2007 659
rect 1435 87 1452 611
rect 2038 87 2055 611
rect 1483 39 2007 56
rect 2181 642 2705 659
rect 2133 87 2150 611
rect 2736 87 2753 611
rect 2181 39 2705 56
rect 2879 642 3403 659
rect 2831 87 2848 611
rect 3434 87 3451 611
rect 2879 39 3403 56
rect 3577 642 4101 659
rect 3529 87 3546 611
rect 4132 87 4149 611
rect 3577 39 4101 56
rect 4275 642 4799 659
rect 4227 87 4244 611
rect 4830 87 4847 611
rect 4275 39 4799 56
rect 4973 642 5497 659
rect 4925 87 4942 611
rect 5528 87 5545 611
rect 4973 39 5497 56
rect 5671 642 6195 659
rect 5623 87 5640 611
rect 6226 87 6243 611
rect 5671 39 6195 56
rect 6369 642 6893 659
rect 6321 87 6338 611
rect 6924 87 6941 611
rect 6369 39 6893 56
rect 7067 642 7591 659
rect 7019 87 7036 611
rect 7622 87 7639 611
rect 7067 39 7591 56
rect 7765 642 8289 659
rect 7717 87 7734 611
rect 8320 87 8337 611
rect 7765 39 8289 56
rect 8463 642 8987 659
rect 8415 87 8432 611
rect 9018 87 9035 611
rect 8463 39 8987 56
rect 9161 642 9685 659
rect 9113 87 9130 611
rect 9716 87 9733 611
rect 9161 39 9685 56
rect 9859 642 10383 659
rect 9811 87 9828 611
rect 10414 87 10431 611
rect 9859 39 10383 56
rect -10383 -56 -9859 -39
rect -10431 -611 -10414 -87
rect -9828 -611 -9811 -87
rect -10383 -659 -9859 -642
rect -9685 -56 -9161 -39
rect -9733 -611 -9716 -87
rect -9130 -611 -9113 -87
rect -9685 -659 -9161 -642
rect -8987 -56 -8463 -39
rect -9035 -611 -9018 -87
rect -8432 -611 -8415 -87
rect -8987 -659 -8463 -642
rect -8289 -56 -7765 -39
rect -8337 -611 -8320 -87
rect -7734 -611 -7717 -87
rect -8289 -659 -7765 -642
rect -7591 -56 -7067 -39
rect -7639 -611 -7622 -87
rect -7036 -611 -7019 -87
rect -7591 -659 -7067 -642
rect -6893 -56 -6369 -39
rect -6941 -611 -6924 -87
rect -6338 -611 -6321 -87
rect -6893 -659 -6369 -642
rect -6195 -56 -5671 -39
rect -6243 -611 -6226 -87
rect -5640 -611 -5623 -87
rect -6195 -659 -5671 -642
rect -5497 -56 -4973 -39
rect -5545 -611 -5528 -87
rect -4942 -611 -4925 -87
rect -5497 -659 -4973 -642
rect -4799 -56 -4275 -39
rect -4847 -611 -4830 -87
rect -4244 -611 -4227 -87
rect -4799 -659 -4275 -642
rect -4101 -56 -3577 -39
rect -4149 -611 -4132 -87
rect -3546 -611 -3529 -87
rect -4101 -659 -3577 -642
rect -3403 -56 -2879 -39
rect -3451 -611 -3434 -87
rect -2848 -611 -2831 -87
rect -3403 -659 -2879 -642
rect -2705 -56 -2181 -39
rect -2753 -611 -2736 -87
rect -2150 -611 -2133 -87
rect -2705 -659 -2181 -642
rect -2007 -56 -1483 -39
rect -2055 -611 -2038 -87
rect -1452 -611 -1435 -87
rect -2007 -659 -1483 -642
rect -1309 -56 -785 -39
rect -1357 -611 -1340 -87
rect -754 -611 -737 -87
rect -1309 -659 -785 -642
rect -611 -56 -87 -39
rect -659 -611 -642 -87
rect -56 -611 -39 -87
rect -611 -659 -87 -642
rect 87 -56 611 -39
rect 39 -611 56 -87
rect 642 -611 659 -87
rect 87 -659 611 -642
rect 785 -56 1309 -39
rect 737 -611 754 -87
rect 1340 -611 1357 -87
rect 785 -659 1309 -642
rect 1483 -56 2007 -39
rect 1435 -611 1452 -87
rect 2038 -611 2055 -87
rect 1483 -659 2007 -642
rect 2181 -56 2705 -39
rect 2133 -611 2150 -87
rect 2736 -611 2753 -87
rect 2181 -659 2705 -642
rect 2879 -56 3403 -39
rect 2831 -611 2848 -87
rect 3434 -611 3451 -87
rect 2879 -659 3403 -642
rect 3577 -56 4101 -39
rect 3529 -611 3546 -87
rect 4132 -611 4149 -87
rect 3577 -659 4101 -642
rect 4275 -56 4799 -39
rect 4227 -611 4244 -87
rect 4830 -611 4847 -87
rect 4275 -659 4799 -642
rect 4973 -56 5497 -39
rect 4925 -611 4942 -87
rect 5528 -611 5545 -87
rect 4973 -659 5497 -642
rect 5671 -56 6195 -39
rect 5623 -611 5640 -87
rect 6226 -611 6243 -87
rect 5671 -659 6195 -642
rect 6369 -56 6893 -39
rect 6321 -611 6338 -87
rect 6924 -611 6941 -87
rect 6369 -659 6893 -642
rect 7067 -56 7591 -39
rect 7019 -611 7036 -87
rect 7622 -611 7639 -87
rect 7067 -659 7591 -642
rect 7765 -56 8289 -39
rect 7717 -611 7734 -87
rect 8320 -611 8337 -87
rect 7765 -659 8289 -642
rect 8463 -56 8987 -39
rect 8415 -611 8432 -87
rect 9018 -611 9035 -87
rect 8463 -659 8987 -642
rect 9161 -56 9685 -39
rect 9113 -611 9130 -87
rect 9716 -611 9733 -87
rect 9161 -659 9685 -642
rect 9859 -56 10383 -39
rect 9811 -611 9828 -87
rect 10414 -611 10431 -87
rect 9859 -659 10383 -642
<< mvpdiode >>
rect -10371 593 -9871 599
rect -10371 105 -10365 593
rect -9877 105 -9871 593
rect -10371 99 -9871 105
rect -9673 593 -9173 599
rect -9673 105 -9667 593
rect -9179 105 -9173 593
rect -9673 99 -9173 105
rect -8975 593 -8475 599
rect -8975 105 -8969 593
rect -8481 105 -8475 593
rect -8975 99 -8475 105
rect -8277 593 -7777 599
rect -8277 105 -8271 593
rect -7783 105 -7777 593
rect -8277 99 -7777 105
rect -7579 593 -7079 599
rect -7579 105 -7573 593
rect -7085 105 -7079 593
rect -7579 99 -7079 105
rect -6881 593 -6381 599
rect -6881 105 -6875 593
rect -6387 105 -6381 593
rect -6881 99 -6381 105
rect -6183 593 -5683 599
rect -6183 105 -6177 593
rect -5689 105 -5683 593
rect -6183 99 -5683 105
rect -5485 593 -4985 599
rect -5485 105 -5479 593
rect -4991 105 -4985 593
rect -5485 99 -4985 105
rect -4787 593 -4287 599
rect -4787 105 -4781 593
rect -4293 105 -4287 593
rect -4787 99 -4287 105
rect -4089 593 -3589 599
rect -4089 105 -4083 593
rect -3595 105 -3589 593
rect -4089 99 -3589 105
rect -3391 593 -2891 599
rect -3391 105 -3385 593
rect -2897 105 -2891 593
rect -3391 99 -2891 105
rect -2693 593 -2193 599
rect -2693 105 -2687 593
rect -2199 105 -2193 593
rect -2693 99 -2193 105
rect -1995 593 -1495 599
rect -1995 105 -1989 593
rect -1501 105 -1495 593
rect -1995 99 -1495 105
rect -1297 593 -797 599
rect -1297 105 -1291 593
rect -803 105 -797 593
rect -1297 99 -797 105
rect -599 593 -99 599
rect -599 105 -593 593
rect -105 105 -99 593
rect -599 99 -99 105
rect 99 593 599 599
rect 99 105 105 593
rect 593 105 599 593
rect 99 99 599 105
rect 797 593 1297 599
rect 797 105 803 593
rect 1291 105 1297 593
rect 797 99 1297 105
rect 1495 593 1995 599
rect 1495 105 1501 593
rect 1989 105 1995 593
rect 1495 99 1995 105
rect 2193 593 2693 599
rect 2193 105 2199 593
rect 2687 105 2693 593
rect 2193 99 2693 105
rect 2891 593 3391 599
rect 2891 105 2897 593
rect 3385 105 3391 593
rect 2891 99 3391 105
rect 3589 593 4089 599
rect 3589 105 3595 593
rect 4083 105 4089 593
rect 3589 99 4089 105
rect 4287 593 4787 599
rect 4287 105 4293 593
rect 4781 105 4787 593
rect 4287 99 4787 105
rect 4985 593 5485 599
rect 4985 105 4991 593
rect 5479 105 5485 593
rect 4985 99 5485 105
rect 5683 593 6183 599
rect 5683 105 5689 593
rect 6177 105 6183 593
rect 5683 99 6183 105
rect 6381 593 6881 599
rect 6381 105 6387 593
rect 6875 105 6881 593
rect 6381 99 6881 105
rect 7079 593 7579 599
rect 7079 105 7085 593
rect 7573 105 7579 593
rect 7079 99 7579 105
rect 7777 593 8277 599
rect 7777 105 7783 593
rect 8271 105 8277 593
rect 7777 99 8277 105
rect 8475 593 8975 599
rect 8475 105 8481 593
rect 8969 105 8975 593
rect 8475 99 8975 105
rect 9173 593 9673 599
rect 9173 105 9179 593
rect 9667 105 9673 593
rect 9173 99 9673 105
rect 9871 593 10371 599
rect 9871 105 9877 593
rect 10365 105 10371 593
rect 9871 99 10371 105
rect -10371 -105 -9871 -99
rect -10371 -593 -10365 -105
rect -9877 -593 -9871 -105
rect -10371 -599 -9871 -593
rect -9673 -105 -9173 -99
rect -9673 -593 -9667 -105
rect -9179 -593 -9173 -105
rect -9673 -599 -9173 -593
rect -8975 -105 -8475 -99
rect -8975 -593 -8969 -105
rect -8481 -593 -8475 -105
rect -8975 -599 -8475 -593
rect -8277 -105 -7777 -99
rect -8277 -593 -8271 -105
rect -7783 -593 -7777 -105
rect -8277 -599 -7777 -593
rect -7579 -105 -7079 -99
rect -7579 -593 -7573 -105
rect -7085 -593 -7079 -105
rect -7579 -599 -7079 -593
rect -6881 -105 -6381 -99
rect -6881 -593 -6875 -105
rect -6387 -593 -6381 -105
rect -6881 -599 -6381 -593
rect -6183 -105 -5683 -99
rect -6183 -593 -6177 -105
rect -5689 -593 -5683 -105
rect -6183 -599 -5683 -593
rect -5485 -105 -4985 -99
rect -5485 -593 -5479 -105
rect -4991 -593 -4985 -105
rect -5485 -599 -4985 -593
rect -4787 -105 -4287 -99
rect -4787 -593 -4781 -105
rect -4293 -593 -4287 -105
rect -4787 -599 -4287 -593
rect -4089 -105 -3589 -99
rect -4089 -593 -4083 -105
rect -3595 -593 -3589 -105
rect -4089 -599 -3589 -593
rect -3391 -105 -2891 -99
rect -3391 -593 -3385 -105
rect -2897 -593 -2891 -105
rect -3391 -599 -2891 -593
rect -2693 -105 -2193 -99
rect -2693 -593 -2687 -105
rect -2199 -593 -2193 -105
rect -2693 -599 -2193 -593
rect -1995 -105 -1495 -99
rect -1995 -593 -1989 -105
rect -1501 -593 -1495 -105
rect -1995 -599 -1495 -593
rect -1297 -105 -797 -99
rect -1297 -593 -1291 -105
rect -803 -593 -797 -105
rect -1297 -599 -797 -593
rect -599 -105 -99 -99
rect -599 -593 -593 -105
rect -105 -593 -99 -105
rect -599 -599 -99 -593
rect 99 -105 599 -99
rect 99 -593 105 -105
rect 593 -593 599 -105
rect 99 -599 599 -593
rect 797 -105 1297 -99
rect 797 -593 803 -105
rect 1291 -593 1297 -105
rect 797 -599 1297 -593
rect 1495 -105 1995 -99
rect 1495 -593 1501 -105
rect 1989 -593 1995 -105
rect 1495 -599 1995 -593
rect 2193 -105 2693 -99
rect 2193 -593 2199 -105
rect 2687 -593 2693 -105
rect 2193 -599 2693 -593
rect 2891 -105 3391 -99
rect 2891 -593 2897 -105
rect 3385 -593 3391 -105
rect 2891 -599 3391 -593
rect 3589 -105 4089 -99
rect 3589 -593 3595 -105
rect 4083 -593 4089 -105
rect 3589 -599 4089 -593
rect 4287 -105 4787 -99
rect 4287 -593 4293 -105
rect 4781 -593 4787 -105
rect 4287 -599 4787 -593
rect 4985 -105 5485 -99
rect 4985 -593 4991 -105
rect 5479 -593 5485 -105
rect 4985 -599 5485 -593
rect 5683 -105 6183 -99
rect 5683 -593 5689 -105
rect 6177 -593 6183 -105
rect 5683 -599 6183 -593
rect 6381 -105 6881 -99
rect 6381 -593 6387 -105
rect 6875 -593 6881 -105
rect 6381 -599 6881 -593
rect 7079 -105 7579 -99
rect 7079 -593 7085 -105
rect 7573 -593 7579 -105
rect 7079 -599 7579 -593
rect 7777 -105 8277 -99
rect 7777 -593 7783 -105
rect 8271 -593 8277 -105
rect 7777 -599 8277 -593
rect 8475 -105 8975 -99
rect 8475 -593 8481 -105
rect 8969 -593 8975 -105
rect 8475 -599 8975 -593
rect 9173 -105 9673 -99
rect 9173 -593 9179 -105
rect 9667 -593 9673 -105
rect 9173 -599 9673 -593
rect 9871 -105 10371 -99
rect 9871 -593 9877 -105
rect 10365 -593 10371 -105
rect 9871 -599 10371 -593
<< mvpdiodec >>
rect -10365 105 -9877 593
rect -9667 105 -9179 593
rect -8969 105 -8481 593
rect -8271 105 -7783 593
rect -7573 105 -7085 593
rect -6875 105 -6387 593
rect -6177 105 -5689 593
rect -5479 105 -4991 593
rect -4781 105 -4293 593
rect -4083 105 -3595 593
rect -3385 105 -2897 593
rect -2687 105 -2199 593
rect -1989 105 -1501 593
rect -1291 105 -803 593
rect -593 105 -105 593
rect 105 105 593 593
rect 803 105 1291 593
rect 1501 105 1989 593
rect 2199 105 2687 593
rect 2897 105 3385 593
rect 3595 105 4083 593
rect 4293 105 4781 593
rect 4991 105 5479 593
rect 5689 105 6177 593
rect 6387 105 6875 593
rect 7085 105 7573 593
rect 7783 105 8271 593
rect 8481 105 8969 593
rect 9179 105 9667 593
rect 9877 105 10365 593
rect -10365 -593 -9877 -105
rect -9667 -593 -9179 -105
rect -8969 -593 -8481 -105
rect -8271 -593 -7783 -105
rect -7573 -593 -7085 -105
rect -6875 -593 -6387 -105
rect -6177 -593 -5689 -105
rect -5479 -593 -4991 -105
rect -4781 -593 -4293 -105
rect -4083 -593 -3595 -105
rect -3385 -593 -2897 -105
rect -2687 -593 -2199 -105
rect -1989 -593 -1501 -105
rect -1291 -593 -803 -105
rect -593 -593 -105 -105
rect 105 -593 593 -105
rect 803 -593 1291 -105
rect 1501 -593 1989 -105
rect 2199 -593 2687 -105
rect 2897 -593 3385 -105
rect 3595 -593 4083 -105
rect 4293 -593 4781 -105
rect 4991 -593 5479 -105
rect 5689 -593 6177 -105
rect 6387 -593 6875 -105
rect 7085 -593 7573 -105
rect 7783 -593 8271 -105
rect 8481 -593 8969 -105
rect 9179 -593 9667 -105
rect 9877 -593 10365 -105
<< locali >>
rect -10536 747 -10488 764
rect 10488 747 10536 764
rect -10536 716 -10519 747
rect 10519 716 10536 747
rect -10431 642 -10383 659
rect -9859 642 -9811 659
rect -10431 611 -10414 642
rect -9828 611 -9811 642
rect -10373 105 -10365 593
rect -9877 105 -9869 593
rect -10431 56 -10414 87
rect -9828 56 -9811 87
rect -10431 39 -10383 56
rect -9859 39 -9811 56
rect -9733 642 -9685 659
rect -9161 642 -9113 659
rect -9733 611 -9716 642
rect -9130 611 -9113 642
rect -9675 105 -9667 593
rect -9179 105 -9171 593
rect -9733 56 -9716 87
rect -9130 56 -9113 87
rect -9733 39 -9685 56
rect -9161 39 -9113 56
rect -9035 642 -8987 659
rect -8463 642 -8415 659
rect -9035 611 -9018 642
rect -8432 611 -8415 642
rect -8977 105 -8969 593
rect -8481 105 -8473 593
rect -9035 56 -9018 87
rect -8432 56 -8415 87
rect -9035 39 -8987 56
rect -8463 39 -8415 56
rect -8337 642 -8289 659
rect -7765 642 -7717 659
rect -8337 611 -8320 642
rect -7734 611 -7717 642
rect -8279 105 -8271 593
rect -7783 105 -7775 593
rect -8337 56 -8320 87
rect -7734 56 -7717 87
rect -8337 39 -8289 56
rect -7765 39 -7717 56
rect -7639 642 -7591 659
rect -7067 642 -7019 659
rect -7639 611 -7622 642
rect -7036 611 -7019 642
rect -7581 105 -7573 593
rect -7085 105 -7077 593
rect -7639 56 -7622 87
rect -7036 56 -7019 87
rect -7639 39 -7591 56
rect -7067 39 -7019 56
rect -6941 642 -6893 659
rect -6369 642 -6321 659
rect -6941 611 -6924 642
rect -6338 611 -6321 642
rect -6883 105 -6875 593
rect -6387 105 -6379 593
rect -6941 56 -6924 87
rect -6338 56 -6321 87
rect -6941 39 -6893 56
rect -6369 39 -6321 56
rect -6243 642 -6195 659
rect -5671 642 -5623 659
rect -6243 611 -6226 642
rect -5640 611 -5623 642
rect -6185 105 -6177 593
rect -5689 105 -5681 593
rect -6243 56 -6226 87
rect -5640 56 -5623 87
rect -6243 39 -6195 56
rect -5671 39 -5623 56
rect -5545 642 -5497 659
rect -4973 642 -4925 659
rect -5545 611 -5528 642
rect -4942 611 -4925 642
rect -5487 105 -5479 593
rect -4991 105 -4983 593
rect -5545 56 -5528 87
rect -4942 56 -4925 87
rect -5545 39 -5497 56
rect -4973 39 -4925 56
rect -4847 642 -4799 659
rect -4275 642 -4227 659
rect -4847 611 -4830 642
rect -4244 611 -4227 642
rect -4789 105 -4781 593
rect -4293 105 -4285 593
rect -4847 56 -4830 87
rect -4244 56 -4227 87
rect -4847 39 -4799 56
rect -4275 39 -4227 56
rect -4149 642 -4101 659
rect -3577 642 -3529 659
rect -4149 611 -4132 642
rect -3546 611 -3529 642
rect -4091 105 -4083 593
rect -3595 105 -3587 593
rect -4149 56 -4132 87
rect -3546 56 -3529 87
rect -4149 39 -4101 56
rect -3577 39 -3529 56
rect -3451 642 -3403 659
rect -2879 642 -2831 659
rect -3451 611 -3434 642
rect -2848 611 -2831 642
rect -3393 105 -3385 593
rect -2897 105 -2889 593
rect -3451 56 -3434 87
rect -2848 56 -2831 87
rect -3451 39 -3403 56
rect -2879 39 -2831 56
rect -2753 642 -2705 659
rect -2181 642 -2133 659
rect -2753 611 -2736 642
rect -2150 611 -2133 642
rect -2695 105 -2687 593
rect -2199 105 -2191 593
rect -2753 56 -2736 87
rect -2150 56 -2133 87
rect -2753 39 -2705 56
rect -2181 39 -2133 56
rect -2055 642 -2007 659
rect -1483 642 -1435 659
rect -2055 611 -2038 642
rect -1452 611 -1435 642
rect -1997 105 -1989 593
rect -1501 105 -1493 593
rect -2055 56 -2038 87
rect -1452 56 -1435 87
rect -2055 39 -2007 56
rect -1483 39 -1435 56
rect -1357 642 -1309 659
rect -785 642 -737 659
rect -1357 611 -1340 642
rect -754 611 -737 642
rect -1299 105 -1291 593
rect -803 105 -795 593
rect -1357 56 -1340 87
rect -754 56 -737 87
rect -1357 39 -1309 56
rect -785 39 -737 56
rect -659 642 -611 659
rect -87 642 -39 659
rect -659 611 -642 642
rect -56 611 -39 642
rect -601 105 -593 593
rect -105 105 -97 593
rect -659 56 -642 87
rect -56 56 -39 87
rect -659 39 -611 56
rect -87 39 -39 56
rect 39 642 87 659
rect 611 642 659 659
rect 39 611 56 642
rect 642 611 659 642
rect 97 105 105 593
rect 593 105 601 593
rect 39 56 56 87
rect 642 56 659 87
rect 39 39 87 56
rect 611 39 659 56
rect 737 642 785 659
rect 1309 642 1357 659
rect 737 611 754 642
rect 1340 611 1357 642
rect 795 105 803 593
rect 1291 105 1299 593
rect 737 56 754 87
rect 1340 56 1357 87
rect 737 39 785 56
rect 1309 39 1357 56
rect 1435 642 1483 659
rect 2007 642 2055 659
rect 1435 611 1452 642
rect 2038 611 2055 642
rect 1493 105 1501 593
rect 1989 105 1997 593
rect 1435 56 1452 87
rect 2038 56 2055 87
rect 1435 39 1483 56
rect 2007 39 2055 56
rect 2133 642 2181 659
rect 2705 642 2753 659
rect 2133 611 2150 642
rect 2736 611 2753 642
rect 2191 105 2199 593
rect 2687 105 2695 593
rect 2133 56 2150 87
rect 2736 56 2753 87
rect 2133 39 2181 56
rect 2705 39 2753 56
rect 2831 642 2879 659
rect 3403 642 3451 659
rect 2831 611 2848 642
rect 3434 611 3451 642
rect 2889 105 2897 593
rect 3385 105 3393 593
rect 2831 56 2848 87
rect 3434 56 3451 87
rect 2831 39 2879 56
rect 3403 39 3451 56
rect 3529 642 3577 659
rect 4101 642 4149 659
rect 3529 611 3546 642
rect 4132 611 4149 642
rect 3587 105 3595 593
rect 4083 105 4091 593
rect 3529 56 3546 87
rect 4132 56 4149 87
rect 3529 39 3577 56
rect 4101 39 4149 56
rect 4227 642 4275 659
rect 4799 642 4847 659
rect 4227 611 4244 642
rect 4830 611 4847 642
rect 4285 105 4293 593
rect 4781 105 4789 593
rect 4227 56 4244 87
rect 4830 56 4847 87
rect 4227 39 4275 56
rect 4799 39 4847 56
rect 4925 642 4973 659
rect 5497 642 5545 659
rect 4925 611 4942 642
rect 5528 611 5545 642
rect 4983 105 4991 593
rect 5479 105 5487 593
rect 4925 56 4942 87
rect 5528 56 5545 87
rect 4925 39 4973 56
rect 5497 39 5545 56
rect 5623 642 5671 659
rect 6195 642 6243 659
rect 5623 611 5640 642
rect 6226 611 6243 642
rect 5681 105 5689 593
rect 6177 105 6185 593
rect 5623 56 5640 87
rect 6226 56 6243 87
rect 5623 39 5671 56
rect 6195 39 6243 56
rect 6321 642 6369 659
rect 6893 642 6941 659
rect 6321 611 6338 642
rect 6924 611 6941 642
rect 6379 105 6387 593
rect 6875 105 6883 593
rect 6321 56 6338 87
rect 6924 56 6941 87
rect 6321 39 6369 56
rect 6893 39 6941 56
rect 7019 642 7067 659
rect 7591 642 7639 659
rect 7019 611 7036 642
rect 7622 611 7639 642
rect 7077 105 7085 593
rect 7573 105 7581 593
rect 7019 56 7036 87
rect 7622 56 7639 87
rect 7019 39 7067 56
rect 7591 39 7639 56
rect 7717 642 7765 659
rect 8289 642 8337 659
rect 7717 611 7734 642
rect 8320 611 8337 642
rect 7775 105 7783 593
rect 8271 105 8279 593
rect 7717 56 7734 87
rect 8320 56 8337 87
rect 7717 39 7765 56
rect 8289 39 8337 56
rect 8415 642 8463 659
rect 8987 642 9035 659
rect 8415 611 8432 642
rect 9018 611 9035 642
rect 8473 105 8481 593
rect 8969 105 8977 593
rect 8415 56 8432 87
rect 9018 56 9035 87
rect 8415 39 8463 56
rect 8987 39 9035 56
rect 9113 642 9161 659
rect 9685 642 9733 659
rect 9113 611 9130 642
rect 9716 611 9733 642
rect 9171 105 9179 593
rect 9667 105 9675 593
rect 9113 56 9130 87
rect 9716 56 9733 87
rect 9113 39 9161 56
rect 9685 39 9733 56
rect 9811 642 9859 659
rect 10383 642 10431 659
rect 9811 611 9828 642
rect 10414 611 10431 642
rect 9869 105 9877 593
rect 10365 105 10373 593
rect 9811 56 9828 87
rect 10414 56 10431 87
rect 9811 39 9859 56
rect 10383 39 10431 56
rect -10431 -56 -10383 -39
rect -9859 -56 -9811 -39
rect -10431 -87 -10414 -56
rect -9828 -87 -9811 -56
rect -10373 -593 -10365 -105
rect -9877 -593 -9869 -105
rect -10431 -642 -10414 -611
rect -9828 -642 -9811 -611
rect -10431 -659 -10383 -642
rect -9859 -659 -9811 -642
rect -9733 -56 -9685 -39
rect -9161 -56 -9113 -39
rect -9733 -87 -9716 -56
rect -9130 -87 -9113 -56
rect -9675 -593 -9667 -105
rect -9179 -593 -9171 -105
rect -9733 -642 -9716 -611
rect -9130 -642 -9113 -611
rect -9733 -659 -9685 -642
rect -9161 -659 -9113 -642
rect -9035 -56 -8987 -39
rect -8463 -56 -8415 -39
rect -9035 -87 -9018 -56
rect -8432 -87 -8415 -56
rect -8977 -593 -8969 -105
rect -8481 -593 -8473 -105
rect -9035 -642 -9018 -611
rect -8432 -642 -8415 -611
rect -9035 -659 -8987 -642
rect -8463 -659 -8415 -642
rect -8337 -56 -8289 -39
rect -7765 -56 -7717 -39
rect -8337 -87 -8320 -56
rect -7734 -87 -7717 -56
rect -8279 -593 -8271 -105
rect -7783 -593 -7775 -105
rect -8337 -642 -8320 -611
rect -7734 -642 -7717 -611
rect -8337 -659 -8289 -642
rect -7765 -659 -7717 -642
rect -7639 -56 -7591 -39
rect -7067 -56 -7019 -39
rect -7639 -87 -7622 -56
rect -7036 -87 -7019 -56
rect -7581 -593 -7573 -105
rect -7085 -593 -7077 -105
rect -7639 -642 -7622 -611
rect -7036 -642 -7019 -611
rect -7639 -659 -7591 -642
rect -7067 -659 -7019 -642
rect -6941 -56 -6893 -39
rect -6369 -56 -6321 -39
rect -6941 -87 -6924 -56
rect -6338 -87 -6321 -56
rect -6883 -593 -6875 -105
rect -6387 -593 -6379 -105
rect -6941 -642 -6924 -611
rect -6338 -642 -6321 -611
rect -6941 -659 -6893 -642
rect -6369 -659 -6321 -642
rect -6243 -56 -6195 -39
rect -5671 -56 -5623 -39
rect -6243 -87 -6226 -56
rect -5640 -87 -5623 -56
rect -6185 -593 -6177 -105
rect -5689 -593 -5681 -105
rect -6243 -642 -6226 -611
rect -5640 -642 -5623 -611
rect -6243 -659 -6195 -642
rect -5671 -659 -5623 -642
rect -5545 -56 -5497 -39
rect -4973 -56 -4925 -39
rect -5545 -87 -5528 -56
rect -4942 -87 -4925 -56
rect -5487 -593 -5479 -105
rect -4991 -593 -4983 -105
rect -5545 -642 -5528 -611
rect -4942 -642 -4925 -611
rect -5545 -659 -5497 -642
rect -4973 -659 -4925 -642
rect -4847 -56 -4799 -39
rect -4275 -56 -4227 -39
rect -4847 -87 -4830 -56
rect -4244 -87 -4227 -56
rect -4789 -593 -4781 -105
rect -4293 -593 -4285 -105
rect -4847 -642 -4830 -611
rect -4244 -642 -4227 -611
rect -4847 -659 -4799 -642
rect -4275 -659 -4227 -642
rect -4149 -56 -4101 -39
rect -3577 -56 -3529 -39
rect -4149 -87 -4132 -56
rect -3546 -87 -3529 -56
rect -4091 -593 -4083 -105
rect -3595 -593 -3587 -105
rect -4149 -642 -4132 -611
rect -3546 -642 -3529 -611
rect -4149 -659 -4101 -642
rect -3577 -659 -3529 -642
rect -3451 -56 -3403 -39
rect -2879 -56 -2831 -39
rect -3451 -87 -3434 -56
rect -2848 -87 -2831 -56
rect -3393 -593 -3385 -105
rect -2897 -593 -2889 -105
rect -3451 -642 -3434 -611
rect -2848 -642 -2831 -611
rect -3451 -659 -3403 -642
rect -2879 -659 -2831 -642
rect -2753 -56 -2705 -39
rect -2181 -56 -2133 -39
rect -2753 -87 -2736 -56
rect -2150 -87 -2133 -56
rect -2695 -593 -2687 -105
rect -2199 -593 -2191 -105
rect -2753 -642 -2736 -611
rect -2150 -642 -2133 -611
rect -2753 -659 -2705 -642
rect -2181 -659 -2133 -642
rect -2055 -56 -2007 -39
rect -1483 -56 -1435 -39
rect -2055 -87 -2038 -56
rect -1452 -87 -1435 -56
rect -1997 -593 -1989 -105
rect -1501 -593 -1493 -105
rect -2055 -642 -2038 -611
rect -1452 -642 -1435 -611
rect -2055 -659 -2007 -642
rect -1483 -659 -1435 -642
rect -1357 -56 -1309 -39
rect -785 -56 -737 -39
rect -1357 -87 -1340 -56
rect -754 -87 -737 -56
rect -1299 -593 -1291 -105
rect -803 -593 -795 -105
rect -1357 -642 -1340 -611
rect -754 -642 -737 -611
rect -1357 -659 -1309 -642
rect -785 -659 -737 -642
rect -659 -56 -611 -39
rect -87 -56 -39 -39
rect -659 -87 -642 -56
rect -56 -87 -39 -56
rect -601 -593 -593 -105
rect -105 -593 -97 -105
rect -659 -642 -642 -611
rect -56 -642 -39 -611
rect -659 -659 -611 -642
rect -87 -659 -39 -642
rect 39 -56 87 -39
rect 611 -56 659 -39
rect 39 -87 56 -56
rect 642 -87 659 -56
rect 97 -593 105 -105
rect 593 -593 601 -105
rect 39 -642 56 -611
rect 642 -642 659 -611
rect 39 -659 87 -642
rect 611 -659 659 -642
rect 737 -56 785 -39
rect 1309 -56 1357 -39
rect 737 -87 754 -56
rect 1340 -87 1357 -56
rect 795 -593 803 -105
rect 1291 -593 1299 -105
rect 737 -642 754 -611
rect 1340 -642 1357 -611
rect 737 -659 785 -642
rect 1309 -659 1357 -642
rect 1435 -56 1483 -39
rect 2007 -56 2055 -39
rect 1435 -87 1452 -56
rect 2038 -87 2055 -56
rect 1493 -593 1501 -105
rect 1989 -593 1997 -105
rect 1435 -642 1452 -611
rect 2038 -642 2055 -611
rect 1435 -659 1483 -642
rect 2007 -659 2055 -642
rect 2133 -56 2181 -39
rect 2705 -56 2753 -39
rect 2133 -87 2150 -56
rect 2736 -87 2753 -56
rect 2191 -593 2199 -105
rect 2687 -593 2695 -105
rect 2133 -642 2150 -611
rect 2736 -642 2753 -611
rect 2133 -659 2181 -642
rect 2705 -659 2753 -642
rect 2831 -56 2879 -39
rect 3403 -56 3451 -39
rect 2831 -87 2848 -56
rect 3434 -87 3451 -56
rect 2889 -593 2897 -105
rect 3385 -593 3393 -105
rect 2831 -642 2848 -611
rect 3434 -642 3451 -611
rect 2831 -659 2879 -642
rect 3403 -659 3451 -642
rect 3529 -56 3577 -39
rect 4101 -56 4149 -39
rect 3529 -87 3546 -56
rect 4132 -87 4149 -56
rect 3587 -593 3595 -105
rect 4083 -593 4091 -105
rect 3529 -642 3546 -611
rect 4132 -642 4149 -611
rect 3529 -659 3577 -642
rect 4101 -659 4149 -642
rect 4227 -56 4275 -39
rect 4799 -56 4847 -39
rect 4227 -87 4244 -56
rect 4830 -87 4847 -56
rect 4285 -593 4293 -105
rect 4781 -593 4789 -105
rect 4227 -642 4244 -611
rect 4830 -642 4847 -611
rect 4227 -659 4275 -642
rect 4799 -659 4847 -642
rect 4925 -56 4973 -39
rect 5497 -56 5545 -39
rect 4925 -87 4942 -56
rect 5528 -87 5545 -56
rect 4983 -593 4991 -105
rect 5479 -593 5487 -105
rect 4925 -642 4942 -611
rect 5528 -642 5545 -611
rect 4925 -659 4973 -642
rect 5497 -659 5545 -642
rect 5623 -56 5671 -39
rect 6195 -56 6243 -39
rect 5623 -87 5640 -56
rect 6226 -87 6243 -56
rect 5681 -593 5689 -105
rect 6177 -593 6185 -105
rect 5623 -642 5640 -611
rect 6226 -642 6243 -611
rect 5623 -659 5671 -642
rect 6195 -659 6243 -642
rect 6321 -56 6369 -39
rect 6893 -56 6941 -39
rect 6321 -87 6338 -56
rect 6924 -87 6941 -56
rect 6379 -593 6387 -105
rect 6875 -593 6883 -105
rect 6321 -642 6338 -611
rect 6924 -642 6941 -611
rect 6321 -659 6369 -642
rect 6893 -659 6941 -642
rect 7019 -56 7067 -39
rect 7591 -56 7639 -39
rect 7019 -87 7036 -56
rect 7622 -87 7639 -56
rect 7077 -593 7085 -105
rect 7573 -593 7581 -105
rect 7019 -642 7036 -611
rect 7622 -642 7639 -611
rect 7019 -659 7067 -642
rect 7591 -659 7639 -642
rect 7717 -56 7765 -39
rect 8289 -56 8337 -39
rect 7717 -87 7734 -56
rect 8320 -87 8337 -56
rect 7775 -593 7783 -105
rect 8271 -593 8279 -105
rect 7717 -642 7734 -611
rect 8320 -642 8337 -611
rect 7717 -659 7765 -642
rect 8289 -659 8337 -642
rect 8415 -56 8463 -39
rect 8987 -56 9035 -39
rect 8415 -87 8432 -56
rect 9018 -87 9035 -56
rect 8473 -593 8481 -105
rect 8969 -593 8977 -105
rect 8415 -642 8432 -611
rect 9018 -642 9035 -611
rect 8415 -659 8463 -642
rect 8987 -659 9035 -642
rect 9113 -56 9161 -39
rect 9685 -56 9733 -39
rect 9113 -87 9130 -56
rect 9716 -87 9733 -56
rect 9171 -593 9179 -105
rect 9667 -593 9675 -105
rect 9113 -642 9130 -611
rect 9716 -642 9733 -611
rect 9113 -659 9161 -642
rect 9685 -659 9733 -642
rect 9811 -56 9859 -39
rect 10383 -56 10431 -39
rect 9811 -87 9828 -56
rect 10414 -87 10431 -56
rect 9869 -593 9877 -105
rect 10365 -593 10373 -105
rect 9811 -642 9828 -611
rect 10414 -642 10431 -611
rect 9811 -659 9859 -642
rect 10383 -659 10431 -642
rect -10536 -747 -10519 -716
rect 10519 -747 10536 -716
rect -10536 -764 -10488 -747
rect 10488 -764 10536 -747
<< viali >>
rect -10365 105 -9877 593
rect -9667 105 -9179 593
rect -8969 105 -8481 593
rect -8271 105 -7783 593
rect -7573 105 -7085 593
rect -6875 105 -6387 593
rect -6177 105 -5689 593
rect -5479 105 -4991 593
rect -4781 105 -4293 593
rect -4083 105 -3595 593
rect -3385 105 -2897 593
rect -2687 105 -2199 593
rect -1989 105 -1501 593
rect -1291 105 -803 593
rect -593 105 -105 593
rect 105 105 593 593
rect 803 105 1291 593
rect 1501 105 1989 593
rect 2199 105 2687 593
rect 2897 105 3385 593
rect 3595 105 4083 593
rect 4293 105 4781 593
rect 4991 105 5479 593
rect 5689 105 6177 593
rect 6387 105 6875 593
rect 7085 105 7573 593
rect 7783 105 8271 593
rect 8481 105 8969 593
rect 9179 105 9667 593
rect 9877 105 10365 593
rect -10365 -593 -9877 -105
rect -9667 -593 -9179 -105
rect -8969 -593 -8481 -105
rect -8271 -593 -7783 -105
rect -7573 -593 -7085 -105
rect -6875 -593 -6387 -105
rect -6177 -593 -5689 -105
rect -5479 -593 -4991 -105
rect -4781 -593 -4293 -105
rect -4083 -593 -3595 -105
rect -3385 -593 -2897 -105
rect -2687 -593 -2199 -105
rect -1989 -593 -1501 -105
rect -1291 -593 -803 -105
rect -593 -593 -105 -105
rect 105 -593 593 -105
rect 803 -593 1291 -105
rect 1501 -593 1989 -105
rect 2199 -593 2687 -105
rect 2897 -593 3385 -105
rect 3595 -593 4083 -105
rect 4293 -593 4781 -105
rect 4991 -593 5479 -105
rect 5689 -593 6177 -105
rect 6387 -593 6875 -105
rect 7085 -593 7573 -105
rect 7783 -593 8271 -105
rect 8481 -593 8969 -105
rect 9179 -593 9667 -105
rect 9877 -593 10365 -105
<< metal1 >>
rect -10371 593 -9871 596
rect -10371 105 -10365 593
rect -9877 105 -9871 593
rect -10371 102 -9871 105
rect -9673 593 -9173 596
rect -9673 105 -9667 593
rect -9179 105 -9173 593
rect -9673 102 -9173 105
rect -8975 593 -8475 596
rect -8975 105 -8969 593
rect -8481 105 -8475 593
rect -8975 102 -8475 105
rect -8277 593 -7777 596
rect -8277 105 -8271 593
rect -7783 105 -7777 593
rect -8277 102 -7777 105
rect -7579 593 -7079 596
rect -7579 105 -7573 593
rect -7085 105 -7079 593
rect -7579 102 -7079 105
rect -6881 593 -6381 596
rect -6881 105 -6875 593
rect -6387 105 -6381 593
rect -6881 102 -6381 105
rect -6183 593 -5683 596
rect -6183 105 -6177 593
rect -5689 105 -5683 593
rect -6183 102 -5683 105
rect -5485 593 -4985 596
rect -5485 105 -5479 593
rect -4991 105 -4985 593
rect -5485 102 -4985 105
rect -4787 593 -4287 596
rect -4787 105 -4781 593
rect -4293 105 -4287 593
rect -4787 102 -4287 105
rect -4089 593 -3589 596
rect -4089 105 -4083 593
rect -3595 105 -3589 593
rect -4089 102 -3589 105
rect -3391 593 -2891 596
rect -3391 105 -3385 593
rect -2897 105 -2891 593
rect -3391 102 -2891 105
rect -2693 593 -2193 596
rect -2693 105 -2687 593
rect -2199 105 -2193 593
rect -2693 102 -2193 105
rect -1995 593 -1495 596
rect -1995 105 -1989 593
rect -1501 105 -1495 593
rect -1995 102 -1495 105
rect -1297 593 -797 596
rect -1297 105 -1291 593
rect -803 105 -797 593
rect -1297 102 -797 105
rect -599 593 -99 596
rect -599 105 -593 593
rect -105 105 -99 593
rect -599 102 -99 105
rect 99 593 599 596
rect 99 105 105 593
rect 593 105 599 593
rect 99 102 599 105
rect 797 593 1297 596
rect 797 105 803 593
rect 1291 105 1297 593
rect 797 102 1297 105
rect 1495 593 1995 596
rect 1495 105 1501 593
rect 1989 105 1995 593
rect 1495 102 1995 105
rect 2193 593 2693 596
rect 2193 105 2199 593
rect 2687 105 2693 593
rect 2193 102 2693 105
rect 2891 593 3391 596
rect 2891 105 2897 593
rect 3385 105 3391 593
rect 2891 102 3391 105
rect 3589 593 4089 596
rect 3589 105 3595 593
rect 4083 105 4089 593
rect 3589 102 4089 105
rect 4287 593 4787 596
rect 4287 105 4293 593
rect 4781 105 4787 593
rect 4287 102 4787 105
rect 4985 593 5485 596
rect 4985 105 4991 593
rect 5479 105 5485 593
rect 4985 102 5485 105
rect 5683 593 6183 596
rect 5683 105 5689 593
rect 6177 105 6183 593
rect 5683 102 6183 105
rect 6381 593 6881 596
rect 6381 105 6387 593
rect 6875 105 6881 593
rect 6381 102 6881 105
rect 7079 593 7579 596
rect 7079 105 7085 593
rect 7573 105 7579 593
rect 7079 102 7579 105
rect 7777 593 8277 596
rect 7777 105 7783 593
rect 8271 105 8277 593
rect 7777 102 8277 105
rect 8475 593 8975 596
rect 8475 105 8481 593
rect 8969 105 8975 593
rect 8475 102 8975 105
rect 9173 593 9673 596
rect 9173 105 9179 593
rect 9667 105 9673 593
rect 9173 102 9673 105
rect 9871 593 10371 596
rect 9871 105 9877 593
rect 10365 105 10371 593
rect 9871 102 10371 105
rect -10371 -105 -9871 -102
rect -10371 -593 -10365 -105
rect -9877 -593 -9871 -105
rect -10371 -596 -9871 -593
rect -9673 -105 -9173 -102
rect -9673 -593 -9667 -105
rect -9179 -593 -9173 -105
rect -9673 -596 -9173 -593
rect -8975 -105 -8475 -102
rect -8975 -593 -8969 -105
rect -8481 -593 -8475 -105
rect -8975 -596 -8475 -593
rect -8277 -105 -7777 -102
rect -8277 -593 -8271 -105
rect -7783 -593 -7777 -105
rect -8277 -596 -7777 -593
rect -7579 -105 -7079 -102
rect -7579 -593 -7573 -105
rect -7085 -593 -7079 -105
rect -7579 -596 -7079 -593
rect -6881 -105 -6381 -102
rect -6881 -593 -6875 -105
rect -6387 -593 -6381 -105
rect -6881 -596 -6381 -593
rect -6183 -105 -5683 -102
rect -6183 -593 -6177 -105
rect -5689 -593 -5683 -105
rect -6183 -596 -5683 -593
rect -5485 -105 -4985 -102
rect -5485 -593 -5479 -105
rect -4991 -593 -4985 -105
rect -5485 -596 -4985 -593
rect -4787 -105 -4287 -102
rect -4787 -593 -4781 -105
rect -4293 -593 -4287 -105
rect -4787 -596 -4287 -593
rect -4089 -105 -3589 -102
rect -4089 -593 -4083 -105
rect -3595 -593 -3589 -105
rect -4089 -596 -3589 -593
rect -3391 -105 -2891 -102
rect -3391 -593 -3385 -105
rect -2897 -593 -2891 -105
rect -3391 -596 -2891 -593
rect -2693 -105 -2193 -102
rect -2693 -593 -2687 -105
rect -2199 -593 -2193 -105
rect -2693 -596 -2193 -593
rect -1995 -105 -1495 -102
rect -1995 -593 -1989 -105
rect -1501 -593 -1495 -105
rect -1995 -596 -1495 -593
rect -1297 -105 -797 -102
rect -1297 -593 -1291 -105
rect -803 -593 -797 -105
rect -1297 -596 -797 -593
rect -599 -105 -99 -102
rect -599 -593 -593 -105
rect -105 -593 -99 -105
rect -599 -596 -99 -593
rect 99 -105 599 -102
rect 99 -593 105 -105
rect 593 -593 599 -105
rect 99 -596 599 -593
rect 797 -105 1297 -102
rect 797 -593 803 -105
rect 1291 -593 1297 -105
rect 797 -596 1297 -593
rect 1495 -105 1995 -102
rect 1495 -593 1501 -105
rect 1989 -593 1995 -105
rect 1495 -596 1995 -593
rect 2193 -105 2693 -102
rect 2193 -593 2199 -105
rect 2687 -593 2693 -105
rect 2193 -596 2693 -593
rect 2891 -105 3391 -102
rect 2891 -593 2897 -105
rect 3385 -593 3391 -105
rect 2891 -596 3391 -593
rect 3589 -105 4089 -102
rect 3589 -593 3595 -105
rect 4083 -593 4089 -105
rect 3589 -596 4089 -593
rect 4287 -105 4787 -102
rect 4287 -593 4293 -105
rect 4781 -593 4787 -105
rect 4287 -596 4787 -593
rect 4985 -105 5485 -102
rect 4985 -593 4991 -105
rect 5479 -593 5485 -105
rect 4985 -596 5485 -593
rect 5683 -105 6183 -102
rect 5683 -593 5689 -105
rect 6177 -593 6183 -105
rect 5683 -596 6183 -593
rect 6381 -105 6881 -102
rect 6381 -593 6387 -105
rect 6875 -593 6881 -105
rect 6381 -596 6881 -593
rect 7079 -105 7579 -102
rect 7079 -593 7085 -105
rect 7573 -593 7579 -105
rect 7079 -596 7579 -593
rect 7777 -105 8277 -102
rect 7777 -593 7783 -105
rect 8271 -593 8277 -105
rect 7777 -596 8277 -593
rect 8475 -105 8975 -102
rect 8475 -593 8481 -105
rect 8969 -593 8975 -105
rect 8475 -596 8975 -593
rect 9173 -105 9673 -102
rect 9173 -593 9179 -105
rect 9667 -593 9673 -105
rect 9173 -596 9673 -593
rect 9871 -105 10371 -102
rect 9871 -593 9877 -105
rect 10365 -593 10371 -105
rect 9871 -596 10371 -593
<< properties >>
string FIXED_BBOX 9819 47 10422 650
string gencell sky130_fd_pr__diode_pd2nw_11v0
string library sky130
string parameters w 5 l 5 area 25.0 peri 20.0 nx 30 ny 2 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 0 compatible {sky130_fd_pr__diode_pd2nw_05v5 sky130_fd_pr__diode_pd2nw_05v5_lvt  sky130_fd_pr__diode_pd2nw_05v5_hvt sky130_fd_pr__diode_pd2nw_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
