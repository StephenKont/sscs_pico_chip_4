magic
tech sky130A
magscale 1 2
timestamp 1666524637
<< error_p >>
rect -70 2800 -10 8200
rect 10 2800 70 8200
rect -70 -2700 -10 2700
rect 10 -2700 70 2700
rect -70 -8200 -10 -2800
rect 10 -8200 70 -2800
<< metal3 >>
rect -5509 8172 -10 8200
rect -5509 2828 -94 8172
rect -30 2828 -10 8172
rect -5509 2800 -10 2828
rect 10 8172 5509 8200
rect 10 2828 5425 8172
rect 5489 2828 5509 8172
rect 10 2800 5509 2828
rect -5509 2672 -10 2700
rect -5509 -2672 -94 2672
rect -30 -2672 -10 2672
rect -5509 -2700 -10 -2672
rect 10 2672 5509 2700
rect 10 -2672 5425 2672
rect 5489 -2672 5509 2672
rect 10 -2700 5509 -2672
rect -5509 -2828 -10 -2800
rect -5509 -8172 -94 -2828
rect -30 -8172 -10 -2828
rect -5509 -8200 -10 -8172
rect 10 -2828 5509 -2800
rect 10 -8172 5425 -2828
rect 5489 -8172 5509 -2828
rect 10 -8200 5509 -8172
<< via3 >>
rect -94 2828 -30 8172
rect 5425 2828 5489 8172
rect -94 -2672 -30 2672
rect 5425 -2672 5489 2672
rect -94 -8172 -30 -2828
rect 5425 -8172 5489 -2828
<< mimcap >>
rect -5409 8060 -209 8100
rect -5409 2940 -5369 8060
rect -249 2940 -209 8060
rect -5409 2900 -209 2940
rect 110 8060 5310 8100
rect 110 2940 150 8060
rect 5270 2940 5310 8060
rect 110 2900 5310 2940
rect -5409 2560 -209 2600
rect -5409 -2560 -5369 2560
rect -249 -2560 -209 2560
rect -5409 -2600 -209 -2560
rect 110 2560 5310 2600
rect 110 -2560 150 2560
rect 5270 -2560 5310 2560
rect 110 -2600 5310 -2560
rect -5409 -2940 -209 -2900
rect -5409 -8060 -5369 -2940
rect -249 -8060 -209 -2940
rect -5409 -8100 -209 -8060
rect 110 -2940 5310 -2900
rect 110 -8060 150 -2940
rect 5270 -8060 5310 -2940
rect 110 -8100 5310 -8060
<< mimcapcontact >>
rect -5369 2940 -249 8060
rect 150 2940 5270 8060
rect -5369 -2560 -249 2560
rect 150 -2560 5270 2560
rect -5369 -8060 -249 -2940
rect 150 -8060 5270 -2940
<< metal4 >>
rect -2861 8061 -2757 8250
rect -141 8188 -37 8250
rect -141 8172 -14 8188
rect -5370 8060 -248 8061
rect -5370 2940 -5369 8060
rect -249 2940 -248 8060
rect -5370 2939 -248 2940
rect -2861 2561 -2757 2939
rect -141 2828 -94 8172
rect -30 2828 -14 8172
rect 2658 8061 2762 8250
rect 5378 8188 5482 8250
rect 5378 8172 5505 8188
rect 149 8060 5271 8061
rect 149 2940 150 8060
rect 5270 2940 5271 8060
rect 149 2939 5271 2940
rect -141 2812 -14 2828
rect -141 2688 -37 2812
rect -141 2672 -14 2688
rect -5370 2560 -248 2561
rect -5370 -2560 -5369 2560
rect -249 -2560 -248 2560
rect -5370 -2561 -248 -2560
rect -2861 -2939 -2757 -2561
rect -141 -2672 -94 2672
rect -30 -2672 -14 2672
rect 2658 2561 2762 2939
rect 5378 2828 5425 8172
rect 5489 2828 5505 8172
rect 5378 2812 5505 2828
rect 5378 2688 5482 2812
rect 5378 2672 5505 2688
rect 149 2560 5271 2561
rect 149 -2560 150 2560
rect 5270 -2560 5271 2560
rect 149 -2561 5271 -2560
rect -141 -2688 -14 -2672
rect -141 -2812 -37 -2688
rect -141 -2828 -14 -2812
rect -5370 -2940 -248 -2939
rect -5370 -8060 -5369 -2940
rect -249 -8060 -248 -2940
rect -5370 -8061 -248 -8060
rect -2861 -8250 -2757 -8061
rect -141 -8172 -94 -2828
rect -30 -8172 -14 -2828
rect 2658 -2939 2762 -2561
rect 5378 -2672 5425 2672
rect 5489 -2672 5505 2672
rect 5378 -2688 5505 -2672
rect 5378 -2812 5482 -2688
rect 5378 -2828 5505 -2812
rect 149 -2940 5271 -2939
rect 149 -8060 150 -2940
rect 5270 -8060 5271 -2940
rect 149 -8061 5271 -8060
rect -141 -8188 -14 -8172
rect -141 -8250 -37 -8188
rect 2658 -8250 2762 -8061
rect 5378 -8172 5425 -2828
rect 5489 -8172 5505 -2828
rect 5378 -8188 5505 -8172
rect 5378 -8250 5482 -8188
<< properties >>
string FIXED_BBOX 10 2800 5410 8200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 26.00 l 26.00 val 1.371k carea 2.00 cperi 0.19 nx 2 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
