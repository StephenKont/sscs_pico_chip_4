magic
tech sky130A
magscale 1 2
timestamp 1665678605
<< error_p >>
rect -607 801 -545 807
rect -479 801 -417 807
rect -351 801 -289 807
rect -223 801 -161 807
rect -95 801 -33 807
rect 33 801 95 807
rect 161 801 223 807
rect 289 801 351 807
rect 417 801 479 807
rect 545 801 607 807
rect -607 767 -595 801
rect -479 767 -467 801
rect -351 767 -339 801
rect -223 767 -211 801
rect -95 767 -83 801
rect 33 767 45 801
rect 161 767 173 801
rect 289 767 301 801
rect 417 767 429 801
rect 545 767 557 801
rect -607 761 -545 767
rect -479 761 -417 767
rect -351 761 -289 767
rect -223 761 -161 767
rect -95 761 -33 767
rect 33 761 95 767
rect 161 761 223 767
rect 289 761 351 767
rect 417 761 479 767
rect 545 761 607 767
rect -607 -767 -545 -761
rect -479 -767 -417 -761
rect -351 -767 -289 -761
rect -223 -767 -161 -761
rect -95 -767 -33 -761
rect 33 -767 95 -761
rect 161 -767 223 -761
rect 289 -767 351 -761
rect 417 -767 479 -761
rect 545 -767 607 -761
rect -607 -801 -595 -767
rect -479 -801 -467 -767
rect -351 -801 -339 -767
rect -223 -801 -211 -767
rect -95 -801 -83 -767
rect 33 -801 45 -767
rect 161 -801 173 -767
rect 289 -801 301 -767
rect 417 -801 429 -767
rect 545 -801 557 -767
rect -607 -807 -545 -801
rect -479 -807 -417 -801
rect -351 -807 -289 -801
rect -223 -807 -161 -801
rect -95 -807 -33 -801
rect 33 -807 95 -801
rect 161 -807 223 -801
rect 289 -807 351 -801
rect 417 -807 479 -801
rect 545 -807 607 -801
<< nwell >>
rect -807 -939 807 939
<< pmoslvt >>
rect -611 -720 -541 720
rect -483 -720 -413 720
rect -355 -720 -285 720
rect -227 -720 -157 720
rect -99 -720 -29 720
rect 29 -720 99 720
rect 157 -720 227 720
rect 285 -720 355 720
rect 413 -720 483 720
rect 541 -720 611 720
<< pdiff >>
rect -669 708 -611 720
rect -669 -708 -657 708
rect -623 -708 -611 708
rect -669 -720 -611 -708
rect -541 708 -483 720
rect -541 -708 -529 708
rect -495 -708 -483 708
rect -541 -720 -483 -708
rect -413 708 -355 720
rect -413 -708 -401 708
rect -367 -708 -355 708
rect -413 -720 -355 -708
rect -285 708 -227 720
rect -285 -708 -273 708
rect -239 -708 -227 708
rect -285 -720 -227 -708
rect -157 708 -99 720
rect -157 -708 -145 708
rect -111 -708 -99 708
rect -157 -720 -99 -708
rect -29 708 29 720
rect -29 -708 -17 708
rect 17 -708 29 708
rect -29 -720 29 -708
rect 99 708 157 720
rect 99 -708 111 708
rect 145 -708 157 708
rect 99 -720 157 -708
rect 227 708 285 720
rect 227 -708 239 708
rect 273 -708 285 708
rect 227 -720 285 -708
rect 355 708 413 720
rect 355 -708 367 708
rect 401 -708 413 708
rect 355 -720 413 -708
rect 483 708 541 720
rect 483 -708 495 708
rect 529 -708 541 708
rect 483 -720 541 -708
rect 611 708 669 720
rect 611 -708 623 708
rect 657 -708 669 708
rect 611 -720 669 -708
<< pdiffc >>
rect -657 -708 -623 708
rect -529 -708 -495 708
rect -401 -708 -367 708
rect -273 -708 -239 708
rect -145 -708 -111 708
rect -17 -708 17 708
rect 111 -708 145 708
rect 239 -708 273 708
rect 367 -708 401 708
rect 495 -708 529 708
rect 623 -708 657 708
<< nsubdiff >>
rect -771 869 -675 903
rect 675 869 771 903
rect -771 807 -737 869
rect 737 807 771 869
rect -771 -869 -737 -807
rect 737 -869 771 -807
rect -771 -903 -675 -869
rect 675 -903 771 -869
<< nsubdiffcont >>
rect -675 869 675 903
rect -771 -807 -737 807
rect 737 -807 771 807
rect -675 -903 675 -869
<< poly >>
rect -611 801 -541 817
rect -611 767 -595 801
rect -557 767 -541 801
rect -611 720 -541 767
rect -483 801 -413 817
rect -483 767 -467 801
rect -429 767 -413 801
rect -483 720 -413 767
rect -355 801 -285 817
rect -355 767 -339 801
rect -301 767 -285 801
rect -355 720 -285 767
rect -227 801 -157 817
rect -227 767 -211 801
rect -173 767 -157 801
rect -227 720 -157 767
rect -99 801 -29 817
rect -99 767 -83 801
rect -45 767 -29 801
rect -99 720 -29 767
rect 29 801 99 817
rect 29 767 45 801
rect 83 767 99 801
rect 29 720 99 767
rect 157 801 227 817
rect 157 767 173 801
rect 211 767 227 801
rect 157 720 227 767
rect 285 801 355 817
rect 285 767 301 801
rect 339 767 355 801
rect 285 720 355 767
rect 413 801 483 817
rect 413 767 429 801
rect 467 767 483 801
rect 413 720 483 767
rect 541 801 611 817
rect 541 767 557 801
rect 595 767 611 801
rect 541 720 611 767
rect -611 -767 -541 -720
rect -611 -801 -595 -767
rect -557 -801 -541 -767
rect -611 -817 -541 -801
rect -483 -767 -413 -720
rect -483 -801 -467 -767
rect -429 -801 -413 -767
rect -483 -817 -413 -801
rect -355 -767 -285 -720
rect -355 -801 -339 -767
rect -301 -801 -285 -767
rect -355 -817 -285 -801
rect -227 -767 -157 -720
rect -227 -801 -211 -767
rect -173 -801 -157 -767
rect -227 -817 -157 -801
rect -99 -767 -29 -720
rect -99 -801 -83 -767
rect -45 -801 -29 -767
rect -99 -817 -29 -801
rect 29 -767 99 -720
rect 29 -801 45 -767
rect 83 -801 99 -767
rect 29 -817 99 -801
rect 157 -767 227 -720
rect 157 -801 173 -767
rect 211 -801 227 -767
rect 157 -817 227 -801
rect 285 -767 355 -720
rect 285 -801 301 -767
rect 339 -801 355 -767
rect 285 -817 355 -801
rect 413 -767 483 -720
rect 413 -801 429 -767
rect 467 -801 483 -767
rect 413 -817 483 -801
rect 541 -767 611 -720
rect 541 -801 557 -767
rect 595 -801 611 -767
rect 541 -817 611 -801
<< polycont >>
rect -595 767 -557 801
rect -467 767 -429 801
rect -339 767 -301 801
rect -211 767 -173 801
rect -83 767 -45 801
rect 45 767 83 801
rect 173 767 211 801
rect 301 767 339 801
rect 429 767 467 801
rect 557 767 595 801
rect -595 -801 -557 -767
rect -467 -801 -429 -767
rect -339 -801 -301 -767
rect -211 -801 -173 -767
rect -83 -801 -45 -767
rect 45 -801 83 -767
rect 173 -801 211 -767
rect 301 -801 339 -767
rect 429 -801 467 -767
rect 557 -801 595 -767
<< locali >>
rect -771 869 -675 903
rect 675 869 771 903
rect -771 807 -737 869
rect 737 807 771 869
rect -611 767 -595 801
rect -557 767 -541 801
rect -483 767 -467 801
rect -429 767 -413 801
rect -355 767 -339 801
rect -301 767 -285 801
rect -227 767 -211 801
rect -173 767 -157 801
rect -99 767 -83 801
rect -45 767 -29 801
rect 29 767 45 801
rect 83 767 99 801
rect 157 767 173 801
rect 211 767 227 801
rect 285 767 301 801
rect 339 767 355 801
rect 413 767 429 801
rect 467 767 483 801
rect 541 767 557 801
rect 595 767 611 801
rect -657 708 -623 724
rect -657 -724 -623 -708
rect -529 708 -495 724
rect -529 -724 -495 -708
rect -401 708 -367 724
rect -401 -724 -367 -708
rect -273 708 -239 724
rect -273 -724 -239 -708
rect -145 708 -111 724
rect -145 -724 -111 -708
rect -17 708 17 724
rect -17 -724 17 -708
rect 111 708 145 724
rect 111 -724 145 -708
rect 239 708 273 724
rect 239 -724 273 -708
rect 367 708 401 724
rect 367 -724 401 -708
rect 495 708 529 724
rect 495 -724 529 -708
rect 623 708 657 724
rect 623 -724 657 -708
rect -611 -801 -595 -767
rect -557 -801 -541 -767
rect -483 -801 -467 -767
rect -429 -801 -413 -767
rect -355 -801 -339 -767
rect -301 -801 -285 -767
rect -227 -801 -211 -767
rect -173 -801 -157 -767
rect -99 -801 -83 -767
rect -45 -801 -29 -767
rect 29 -801 45 -767
rect 83 -801 99 -767
rect 157 -801 173 -767
rect 211 -801 227 -767
rect 285 -801 301 -767
rect 339 -801 355 -767
rect 413 -801 429 -767
rect 467 -801 483 -767
rect 541 -801 557 -767
rect 595 -801 611 -767
rect -771 -869 -737 -807
rect 737 -869 771 -807
rect -771 -903 -675 -869
rect 675 -903 771 -869
<< viali >>
rect -595 767 -557 801
rect -467 767 -429 801
rect -339 767 -301 801
rect -211 767 -173 801
rect -83 767 -45 801
rect 45 767 83 801
rect 173 767 211 801
rect 301 767 339 801
rect 429 767 467 801
rect 557 767 595 801
rect -657 -708 -623 708
rect -529 -708 -495 708
rect -401 -708 -367 708
rect -273 -708 -239 708
rect -145 -708 -111 708
rect -17 -708 17 708
rect 111 -708 145 708
rect 239 -708 273 708
rect 367 -708 401 708
rect 495 -708 529 708
rect 623 -708 657 708
rect -595 -801 -557 -767
rect -467 -801 -429 -767
rect -339 -801 -301 -767
rect -211 -801 -173 -767
rect -83 -801 -45 -767
rect 45 -801 83 -767
rect 173 -801 211 -767
rect 301 -801 339 -767
rect 429 -801 467 -767
rect 557 -801 595 -767
<< metal1 >>
rect -607 801 -545 807
rect -607 767 -595 801
rect -557 767 -545 801
rect -607 761 -545 767
rect -479 801 -417 807
rect -479 767 -467 801
rect -429 767 -417 801
rect -479 761 -417 767
rect -351 801 -289 807
rect -351 767 -339 801
rect -301 767 -289 801
rect -351 761 -289 767
rect -223 801 -161 807
rect -223 767 -211 801
rect -173 767 -161 801
rect -223 761 -161 767
rect -95 801 -33 807
rect -95 767 -83 801
rect -45 767 -33 801
rect -95 761 -33 767
rect 33 801 95 807
rect 33 767 45 801
rect 83 767 95 801
rect 33 761 95 767
rect 161 801 223 807
rect 161 767 173 801
rect 211 767 223 801
rect 161 761 223 767
rect 289 801 351 807
rect 289 767 301 801
rect 339 767 351 801
rect 289 761 351 767
rect 417 801 479 807
rect 417 767 429 801
rect 467 767 479 801
rect 417 761 479 767
rect 545 801 607 807
rect 545 767 557 801
rect 595 767 607 801
rect 545 761 607 767
rect -663 708 -617 720
rect -663 -708 -657 708
rect -623 -708 -617 708
rect -663 -720 -617 -708
rect -535 708 -489 720
rect -535 -708 -529 708
rect -495 -708 -489 708
rect -535 -720 -489 -708
rect -407 708 -361 720
rect -407 -708 -401 708
rect -367 -708 -361 708
rect -407 -720 -361 -708
rect -279 708 -233 720
rect -279 -708 -273 708
rect -239 -708 -233 708
rect -279 -720 -233 -708
rect -151 708 -105 720
rect -151 -708 -145 708
rect -111 -708 -105 708
rect -151 -720 -105 -708
rect -23 708 23 720
rect -23 -708 -17 708
rect 17 -708 23 708
rect -23 -720 23 -708
rect 105 708 151 720
rect 105 -708 111 708
rect 145 -708 151 708
rect 105 -720 151 -708
rect 233 708 279 720
rect 233 -708 239 708
rect 273 -708 279 708
rect 233 -720 279 -708
rect 361 708 407 720
rect 361 -708 367 708
rect 401 -708 407 708
rect 361 -720 407 -708
rect 489 708 535 720
rect 489 -708 495 708
rect 529 -708 535 708
rect 489 -720 535 -708
rect 617 708 663 720
rect 617 -708 623 708
rect 657 -708 663 708
rect 617 -720 663 -708
rect -607 -767 -545 -761
rect -607 -801 -595 -767
rect -557 -801 -545 -767
rect -607 -807 -545 -801
rect -479 -767 -417 -761
rect -479 -801 -467 -767
rect -429 -801 -417 -767
rect -479 -807 -417 -801
rect -351 -767 -289 -761
rect -351 -801 -339 -767
rect -301 -801 -289 -767
rect -351 -807 -289 -801
rect -223 -767 -161 -761
rect -223 -801 -211 -767
rect -173 -801 -161 -767
rect -223 -807 -161 -801
rect -95 -767 -33 -761
rect -95 -801 -83 -767
rect -45 -801 -33 -767
rect -95 -807 -33 -801
rect 33 -767 95 -761
rect 33 -801 45 -767
rect 83 -801 95 -767
rect 33 -807 95 -801
rect 161 -767 223 -761
rect 161 -801 173 -767
rect 211 -801 223 -767
rect 161 -807 223 -801
rect 289 -767 351 -761
rect 289 -801 301 -767
rect 339 -801 351 -767
rect 289 -807 351 -801
rect 417 -767 479 -761
rect 417 -801 429 -767
rect 467 -801 479 -767
rect 417 -807 479 -801
rect 545 -767 607 -761
rect 545 -801 557 -767
rect 595 -801 607 -767
rect 545 -807 607 -801
<< properties >>
string FIXED_BBOX -754 -886 754 886
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 7.2 l 0.35 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
