magic
tech sky130A
magscale 1 2
timestamp 1664842101
<< pwell >>
rect -6519 -2478 6519 2478
<< mvnmos >>
rect -6291 1420 -6191 2220
rect -6133 1420 -6033 2220
rect -5975 1420 -5875 2220
rect -5817 1420 -5717 2220
rect -5659 1420 -5559 2220
rect -5501 1420 -5401 2220
rect -5343 1420 -5243 2220
rect -5185 1420 -5085 2220
rect -5027 1420 -4927 2220
rect -4869 1420 -4769 2220
rect -4711 1420 -4611 2220
rect -4553 1420 -4453 2220
rect -4395 1420 -4295 2220
rect -4237 1420 -4137 2220
rect -4079 1420 -3979 2220
rect -3921 1420 -3821 2220
rect -3763 1420 -3663 2220
rect -3605 1420 -3505 2220
rect -3447 1420 -3347 2220
rect -3289 1420 -3189 2220
rect -3131 1420 -3031 2220
rect -2973 1420 -2873 2220
rect -2815 1420 -2715 2220
rect -2657 1420 -2557 2220
rect -2499 1420 -2399 2220
rect -2341 1420 -2241 2220
rect -2183 1420 -2083 2220
rect -2025 1420 -1925 2220
rect -1867 1420 -1767 2220
rect -1709 1420 -1609 2220
rect -1551 1420 -1451 2220
rect -1393 1420 -1293 2220
rect -1235 1420 -1135 2220
rect -1077 1420 -977 2220
rect -919 1420 -819 2220
rect -761 1420 -661 2220
rect -603 1420 -503 2220
rect -445 1420 -345 2220
rect -287 1420 -187 2220
rect -129 1420 -29 2220
rect 29 1420 129 2220
rect 187 1420 287 2220
rect 345 1420 445 2220
rect 503 1420 603 2220
rect 661 1420 761 2220
rect 819 1420 919 2220
rect 977 1420 1077 2220
rect 1135 1420 1235 2220
rect 1293 1420 1393 2220
rect 1451 1420 1551 2220
rect 1609 1420 1709 2220
rect 1767 1420 1867 2220
rect 1925 1420 2025 2220
rect 2083 1420 2183 2220
rect 2241 1420 2341 2220
rect 2399 1420 2499 2220
rect 2557 1420 2657 2220
rect 2715 1420 2815 2220
rect 2873 1420 2973 2220
rect 3031 1420 3131 2220
rect 3189 1420 3289 2220
rect 3347 1420 3447 2220
rect 3505 1420 3605 2220
rect 3663 1420 3763 2220
rect 3821 1420 3921 2220
rect 3979 1420 4079 2220
rect 4137 1420 4237 2220
rect 4295 1420 4395 2220
rect 4453 1420 4553 2220
rect 4611 1420 4711 2220
rect 4769 1420 4869 2220
rect 4927 1420 5027 2220
rect 5085 1420 5185 2220
rect 5243 1420 5343 2220
rect 5401 1420 5501 2220
rect 5559 1420 5659 2220
rect 5717 1420 5817 2220
rect 5875 1420 5975 2220
rect 6033 1420 6133 2220
rect 6191 1420 6291 2220
rect -6291 510 -6191 1310
rect -6133 510 -6033 1310
rect -5975 510 -5875 1310
rect -5817 510 -5717 1310
rect -5659 510 -5559 1310
rect -5501 510 -5401 1310
rect -5343 510 -5243 1310
rect -5185 510 -5085 1310
rect -5027 510 -4927 1310
rect -4869 510 -4769 1310
rect -4711 510 -4611 1310
rect -4553 510 -4453 1310
rect -4395 510 -4295 1310
rect -4237 510 -4137 1310
rect -4079 510 -3979 1310
rect -3921 510 -3821 1310
rect -3763 510 -3663 1310
rect -3605 510 -3505 1310
rect -3447 510 -3347 1310
rect -3289 510 -3189 1310
rect -3131 510 -3031 1310
rect -2973 510 -2873 1310
rect -2815 510 -2715 1310
rect -2657 510 -2557 1310
rect -2499 510 -2399 1310
rect -2341 510 -2241 1310
rect -2183 510 -2083 1310
rect -2025 510 -1925 1310
rect -1867 510 -1767 1310
rect -1709 510 -1609 1310
rect -1551 510 -1451 1310
rect -1393 510 -1293 1310
rect -1235 510 -1135 1310
rect -1077 510 -977 1310
rect -919 510 -819 1310
rect -761 510 -661 1310
rect -603 510 -503 1310
rect -445 510 -345 1310
rect -287 510 -187 1310
rect -129 510 -29 1310
rect 29 510 129 1310
rect 187 510 287 1310
rect 345 510 445 1310
rect 503 510 603 1310
rect 661 510 761 1310
rect 819 510 919 1310
rect 977 510 1077 1310
rect 1135 510 1235 1310
rect 1293 510 1393 1310
rect 1451 510 1551 1310
rect 1609 510 1709 1310
rect 1767 510 1867 1310
rect 1925 510 2025 1310
rect 2083 510 2183 1310
rect 2241 510 2341 1310
rect 2399 510 2499 1310
rect 2557 510 2657 1310
rect 2715 510 2815 1310
rect 2873 510 2973 1310
rect 3031 510 3131 1310
rect 3189 510 3289 1310
rect 3347 510 3447 1310
rect 3505 510 3605 1310
rect 3663 510 3763 1310
rect 3821 510 3921 1310
rect 3979 510 4079 1310
rect 4137 510 4237 1310
rect 4295 510 4395 1310
rect 4453 510 4553 1310
rect 4611 510 4711 1310
rect 4769 510 4869 1310
rect 4927 510 5027 1310
rect 5085 510 5185 1310
rect 5243 510 5343 1310
rect 5401 510 5501 1310
rect 5559 510 5659 1310
rect 5717 510 5817 1310
rect 5875 510 5975 1310
rect 6033 510 6133 1310
rect 6191 510 6291 1310
rect -6291 -400 -6191 400
rect -6133 -400 -6033 400
rect -5975 -400 -5875 400
rect -5817 -400 -5717 400
rect -5659 -400 -5559 400
rect -5501 -400 -5401 400
rect -5343 -400 -5243 400
rect -5185 -400 -5085 400
rect -5027 -400 -4927 400
rect -4869 -400 -4769 400
rect -4711 -400 -4611 400
rect -4553 -400 -4453 400
rect -4395 -400 -4295 400
rect -4237 -400 -4137 400
rect -4079 -400 -3979 400
rect -3921 -400 -3821 400
rect -3763 -400 -3663 400
rect -3605 -400 -3505 400
rect -3447 -400 -3347 400
rect -3289 -400 -3189 400
rect -3131 -400 -3031 400
rect -2973 -400 -2873 400
rect -2815 -400 -2715 400
rect -2657 -400 -2557 400
rect -2499 -400 -2399 400
rect -2341 -400 -2241 400
rect -2183 -400 -2083 400
rect -2025 -400 -1925 400
rect -1867 -400 -1767 400
rect -1709 -400 -1609 400
rect -1551 -400 -1451 400
rect -1393 -400 -1293 400
rect -1235 -400 -1135 400
rect -1077 -400 -977 400
rect -919 -400 -819 400
rect -761 -400 -661 400
rect -603 -400 -503 400
rect -445 -400 -345 400
rect -287 -400 -187 400
rect -129 -400 -29 400
rect 29 -400 129 400
rect 187 -400 287 400
rect 345 -400 445 400
rect 503 -400 603 400
rect 661 -400 761 400
rect 819 -400 919 400
rect 977 -400 1077 400
rect 1135 -400 1235 400
rect 1293 -400 1393 400
rect 1451 -400 1551 400
rect 1609 -400 1709 400
rect 1767 -400 1867 400
rect 1925 -400 2025 400
rect 2083 -400 2183 400
rect 2241 -400 2341 400
rect 2399 -400 2499 400
rect 2557 -400 2657 400
rect 2715 -400 2815 400
rect 2873 -400 2973 400
rect 3031 -400 3131 400
rect 3189 -400 3289 400
rect 3347 -400 3447 400
rect 3505 -400 3605 400
rect 3663 -400 3763 400
rect 3821 -400 3921 400
rect 3979 -400 4079 400
rect 4137 -400 4237 400
rect 4295 -400 4395 400
rect 4453 -400 4553 400
rect 4611 -400 4711 400
rect 4769 -400 4869 400
rect 4927 -400 5027 400
rect 5085 -400 5185 400
rect 5243 -400 5343 400
rect 5401 -400 5501 400
rect 5559 -400 5659 400
rect 5717 -400 5817 400
rect 5875 -400 5975 400
rect 6033 -400 6133 400
rect 6191 -400 6291 400
rect -6291 -1310 -6191 -510
rect -6133 -1310 -6033 -510
rect -5975 -1310 -5875 -510
rect -5817 -1310 -5717 -510
rect -5659 -1310 -5559 -510
rect -5501 -1310 -5401 -510
rect -5343 -1310 -5243 -510
rect -5185 -1310 -5085 -510
rect -5027 -1310 -4927 -510
rect -4869 -1310 -4769 -510
rect -4711 -1310 -4611 -510
rect -4553 -1310 -4453 -510
rect -4395 -1310 -4295 -510
rect -4237 -1310 -4137 -510
rect -4079 -1310 -3979 -510
rect -3921 -1310 -3821 -510
rect -3763 -1310 -3663 -510
rect -3605 -1310 -3505 -510
rect -3447 -1310 -3347 -510
rect -3289 -1310 -3189 -510
rect -3131 -1310 -3031 -510
rect -2973 -1310 -2873 -510
rect -2815 -1310 -2715 -510
rect -2657 -1310 -2557 -510
rect -2499 -1310 -2399 -510
rect -2341 -1310 -2241 -510
rect -2183 -1310 -2083 -510
rect -2025 -1310 -1925 -510
rect -1867 -1310 -1767 -510
rect -1709 -1310 -1609 -510
rect -1551 -1310 -1451 -510
rect -1393 -1310 -1293 -510
rect -1235 -1310 -1135 -510
rect -1077 -1310 -977 -510
rect -919 -1310 -819 -510
rect -761 -1310 -661 -510
rect -603 -1310 -503 -510
rect -445 -1310 -345 -510
rect -287 -1310 -187 -510
rect -129 -1310 -29 -510
rect 29 -1310 129 -510
rect 187 -1310 287 -510
rect 345 -1310 445 -510
rect 503 -1310 603 -510
rect 661 -1310 761 -510
rect 819 -1310 919 -510
rect 977 -1310 1077 -510
rect 1135 -1310 1235 -510
rect 1293 -1310 1393 -510
rect 1451 -1310 1551 -510
rect 1609 -1310 1709 -510
rect 1767 -1310 1867 -510
rect 1925 -1310 2025 -510
rect 2083 -1310 2183 -510
rect 2241 -1310 2341 -510
rect 2399 -1310 2499 -510
rect 2557 -1310 2657 -510
rect 2715 -1310 2815 -510
rect 2873 -1310 2973 -510
rect 3031 -1310 3131 -510
rect 3189 -1310 3289 -510
rect 3347 -1310 3447 -510
rect 3505 -1310 3605 -510
rect 3663 -1310 3763 -510
rect 3821 -1310 3921 -510
rect 3979 -1310 4079 -510
rect 4137 -1310 4237 -510
rect 4295 -1310 4395 -510
rect 4453 -1310 4553 -510
rect 4611 -1310 4711 -510
rect 4769 -1310 4869 -510
rect 4927 -1310 5027 -510
rect 5085 -1310 5185 -510
rect 5243 -1310 5343 -510
rect 5401 -1310 5501 -510
rect 5559 -1310 5659 -510
rect 5717 -1310 5817 -510
rect 5875 -1310 5975 -510
rect 6033 -1310 6133 -510
rect 6191 -1310 6291 -510
rect -6291 -2220 -6191 -1420
rect -6133 -2220 -6033 -1420
rect -5975 -2220 -5875 -1420
rect -5817 -2220 -5717 -1420
rect -5659 -2220 -5559 -1420
rect -5501 -2220 -5401 -1420
rect -5343 -2220 -5243 -1420
rect -5185 -2220 -5085 -1420
rect -5027 -2220 -4927 -1420
rect -4869 -2220 -4769 -1420
rect -4711 -2220 -4611 -1420
rect -4553 -2220 -4453 -1420
rect -4395 -2220 -4295 -1420
rect -4237 -2220 -4137 -1420
rect -4079 -2220 -3979 -1420
rect -3921 -2220 -3821 -1420
rect -3763 -2220 -3663 -1420
rect -3605 -2220 -3505 -1420
rect -3447 -2220 -3347 -1420
rect -3289 -2220 -3189 -1420
rect -3131 -2220 -3031 -1420
rect -2973 -2220 -2873 -1420
rect -2815 -2220 -2715 -1420
rect -2657 -2220 -2557 -1420
rect -2499 -2220 -2399 -1420
rect -2341 -2220 -2241 -1420
rect -2183 -2220 -2083 -1420
rect -2025 -2220 -1925 -1420
rect -1867 -2220 -1767 -1420
rect -1709 -2220 -1609 -1420
rect -1551 -2220 -1451 -1420
rect -1393 -2220 -1293 -1420
rect -1235 -2220 -1135 -1420
rect -1077 -2220 -977 -1420
rect -919 -2220 -819 -1420
rect -761 -2220 -661 -1420
rect -603 -2220 -503 -1420
rect -445 -2220 -345 -1420
rect -287 -2220 -187 -1420
rect -129 -2220 -29 -1420
rect 29 -2220 129 -1420
rect 187 -2220 287 -1420
rect 345 -2220 445 -1420
rect 503 -2220 603 -1420
rect 661 -2220 761 -1420
rect 819 -2220 919 -1420
rect 977 -2220 1077 -1420
rect 1135 -2220 1235 -1420
rect 1293 -2220 1393 -1420
rect 1451 -2220 1551 -1420
rect 1609 -2220 1709 -1420
rect 1767 -2220 1867 -1420
rect 1925 -2220 2025 -1420
rect 2083 -2220 2183 -1420
rect 2241 -2220 2341 -1420
rect 2399 -2220 2499 -1420
rect 2557 -2220 2657 -1420
rect 2715 -2220 2815 -1420
rect 2873 -2220 2973 -1420
rect 3031 -2220 3131 -1420
rect 3189 -2220 3289 -1420
rect 3347 -2220 3447 -1420
rect 3505 -2220 3605 -1420
rect 3663 -2220 3763 -1420
rect 3821 -2220 3921 -1420
rect 3979 -2220 4079 -1420
rect 4137 -2220 4237 -1420
rect 4295 -2220 4395 -1420
rect 4453 -2220 4553 -1420
rect 4611 -2220 4711 -1420
rect 4769 -2220 4869 -1420
rect 4927 -2220 5027 -1420
rect 5085 -2220 5185 -1420
rect 5243 -2220 5343 -1420
rect 5401 -2220 5501 -1420
rect 5559 -2220 5659 -1420
rect 5717 -2220 5817 -1420
rect 5875 -2220 5975 -1420
rect 6033 -2220 6133 -1420
rect 6191 -2220 6291 -1420
<< mvndiff >>
rect -6349 2208 -6291 2220
rect -6349 1432 -6337 2208
rect -6303 1432 -6291 2208
rect -6349 1420 -6291 1432
rect -6191 2208 -6133 2220
rect -6191 1432 -6179 2208
rect -6145 1432 -6133 2208
rect -6191 1420 -6133 1432
rect -6033 2208 -5975 2220
rect -6033 1432 -6021 2208
rect -5987 1432 -5975 2208
rect -6033 1420 -5975 1432
rect -5875 2208 -5817 2220
rect -5875 1432 -5863 2208
rect -5829 1432 -5817 2208
rect -5875 1420 -5817 1432
rect -5717 2208 -5659 2220
rect -5717 1432 -5705 2208
rect -5671 1432 -5659 2208
rect -5717 1420 -5659 1432
rect -5559 2208 -5501 2220
rect -5559 1432 -5547 2208
rect -5513 1432 -5501 2208
rect -5559 1420 -5501 1432
rect -5401 2208 -5343 2220
rect -5401 1432 -5389 2208
rect -5355 1432 -5343 2208
rect -5401 1420 -5343 1432
rect -5243 2208 -5185 2220
rect -5243 1432 -5231 2208
rect -5197 1432 -5185 2208
rect -5243 1420 -5185 1432
rect -5085 2208 -5027 2220
rect -5085 1432 -5073 2208
rect -5039 1432 -5027 2208
rect -5085 1420 -5027 1432
rect -4927 2208 -4869 2220
rect -4927 1432 -4915 2208
rect -4881 1432 -4869 2208
rect -4927 1420 -4869 1432
rect -4769 2208 -4711 2220
rect -4769 1432 -4757 2208
rect -4723 1432 -4711 2208
rect -4769 1420 -4711 1432
rect -4611 2208 -4553 2220
rect -4611 1432 -4599 2208
rect -4565 1432 -4553 2208
rect -4611 1420 -4553 1432
rect -4453 2208 -4395 2220
rect -4453 1432 -4441 2208
rect -4407 1432 -4395 2208
rect -4453 1420 -4395 1432
rect -4295 2208 -4237 2220
rect -4295 1432 -4283 2208
rect -4249 1432 -4237 2208
rect -4295 1420 -4237 1432
rect -4137 2208 -4079 2220
rect -4137 1432 -4125 2208
rect -4091 1432 -4079 2208
rect -4137 1420 -4079 1432
rect -3979 2208 -3921 2220
rect -3979 1432 -3967 2208
rect -3933 1432 -3921 2208
rect -3979 1420 -3921 1432
rect -3821 2208 -3763 2220
rect -3821 1432 -3809 2208
rect -3775 1432 -3763 2208
rect -3821 1420 -3763 1432
rect -3663 2208 -3605 2220
rect -3663 1432 -3651 2208
rect -3617 1432 -3605 2208
rect -3663 1420 -3605 1432
rect -3505 2208 -3447 2220
rect -3505 1432 -3493 2208
rect -3459 1432 -3447 2208
rect -3505 1420 -3447 1432
rect -3347 2208 -3289 2220
rect -3347 1432 -3335 2208
rect -3301 1432 -3289 2208
rect -3347 1420 -3289 1432
rect -3189 2208 -3131 2220
rect -3189 1432 -3177 2208
rect -3143 1432 -3131 2208
rect -3189 1420 -3131 1432
rect -3031 2208 -2973 2220
rect -3031 1432 -3019 2208
rect -2985 1432 -2973 2208
rect -3031 1420 -2973 1432
rect -2873 2208 -2815 2220
rect -2873 1432 -2861 2208
rect -2827 1432 -2815 2208
rect -2873 1420 -2815 1432
rect -2715 2208 -2657 2220
rect -2715 1432 -2703 2208
rect -2669 1432 -2657 2208
rect -2715 1420 -2657 1432
rect -2557 2208 -2499 2220
rect -2557 1432 -2545 2208
rect -2511 1432 -2499 2208
rect -2557 1420 -2499 1432
rect -2399 2208 -2341 2220
rect -2399 1432 -2387 2208
rect -2353 1432 -2341 2208
rect -2399 1420 -2341 1432
rect -2241 2208 -2183 2220
rect -2241 1432 -2229 2208
rect -2195 1432 -2183 2208
rect -2241 1420 -2183 1432
rect -2083 2208 -2025 2220
rect -2083 1432 -2071 2208
rect -2037 1432 -2025 2208
rect -2083 1420 -2025 1432
rect -1925 2208 -1867 2220
rect -1925 1432 -1913 2208
rect -1879 1432 -1867 2208
rect -1925 1420 -1867 1432
rect -1767 2208 -1709 2220
rect -1767 1432 -1755 2208
rect -1721 1432 -1709 2208
rect -1767 1420 -1709 1432
rect -1609 2208 -1551 2220
rect -1609 1432 -1597 2208
rect -1563 1432 -1551 2208
rect -1609 1420 -1551 1432
rect -1451 2208 -1393 2220
rect -1451 1432 -1439 2208
rect -1405 1432 -1393 2208
rect -1451 1420 -1393 1432
rect -1293 2208 -1235 2220
rect -1293 1432 -1281 2208
rect -1247 1432 -1235 2208
rect -1293 1420 -1235 1432
rect -1135 2208 -1077 2220
rect -1135 1432 -1123 2208
rect -1089 1432 -1077 2208
rect -1135 1420 -1077 1432
rect -977 2208 -919 2220
rect -977 1432 -965 2208
rect -931 1432 -919 2208
rect -977 1420 -919 1432
rect -819 2208 -761 2220
rect -819 1432 -807 2208
rect -773 1432 -761 2208
rect -819 1420 -761 1432
rect -661 2208 -603 2220
rect -661 1432 -649 2208
rect -615 1432 -603 2208
rect -661 1420 -603 1432
rect -503 2208 -445 2220
rect -503 1432 -491 2208
rect -457 1432 -445 2208
rect -503 1420 -445 1432
rect -345 2208 -287 2220
rect -345 1432 -333 2208
rect -299 1432 -287 2208
rect -345 1420 -287 1432
rect -187 2208 -129 2220
rect -187 1432 -175 2208
rect -141 1432 -129 2208
rect -187 1420 -129 1432
rect -29 2208 29 2220
rect -29 1432 -17 2208
rect 17 1432 29 2208
rect -29 1420 29 1432
rect 129 2208 187 2220
rect 129 1432 141 2208
rect 175 1432 187 2208
rect 129 1420 187 1432
rect 287 2208 345 2220
rect 287 1432 299 2208
rect 333 1432 345 2208
rect 287 1420 345 1432
rect 445 2208 503 2220
rect 445 1432 457 2208
rect 491 1432 503 2208
rect 445 1420 503 1432
rect 603 2208 661 2220
rect 603 1432 615 2208
rect 649 1432 661 2208
rect 603 1420 661 1432
rect 761 2208 819 2220
rect 761 1432 773 2208
rect 807 1432 819 2208
rect 761 1420 819 1432
rect 919 2208 977 2220
rect 919 1432 931 2208
rect 965 1432 977 2208
rect 919 1420 977 1432
rect 1077 2208 1135 2220
rect 1077 1432 1089 2208
rect 1123 1432 1135 2208
rect 1077 1420 1135 1432
rect 1235 2208 1293 2220
rect 1235 1432 1247 2208
rect 1281 1432 1293 2208
rect 1235 1420 1293 1432
rect 1393 2208 1451 2220
rect 1393 1432 1405 2208
rect 1439 1432 1451 2208
rect 1393 1420 1451 1432
rect 1551 2208 1609 2220
rect 1551 1432 1563 2208
rect 1597 1432 1609 2208
rect 1551 1420 1609 1432
rect 1709 2208 1767 2220
rect 1709 1432 1721 2208
rect 1755 1432 1767 2208
rect 1709 1420 1767 1432
rect 1867 2208 1925 2220
rect 1867 1432 1879 2208
rect 1913 1432 1925 2208
rect 1867 1420 1925 1432
rect 2025 2208 2083 2220
rect 2025 1432 2037 2208
rect 2071 1432 2083 2208
rect 2025 1420 2083 1432
rect 2183 2208 2241 2220
rect 2183 1432 2195 2208
rect 2229 1432 2241 2208
rect 2183 1420 2241 1432
rect 2341 2208 2399 2220
rect 2341 1432 2353 2208
rect 2387 1432 2399 2208
rect 2341 1420 2399 1432
rect 2499 2208 2557 2220
rect 2499 1432 2511 2208
rect 2545 1432 2557 2208
rect 2499 1420 2557 1432
rect 2657 2208 2715 2220
rect 2657 1432 2669 2208
rect 2703 1432 2715 2208
rect 2657 1420 2715 1432
rect 2815 2208 2873 2220
rect 2815 1432 2827 2208
rect 2861 1432 2873 2208
rect 2815 1420 2873 1432
rect 2973 2208 3031 2220
rect 2973 1432 2985 2208
rect 3019 1432 3031 2208
rect 2973 1420 3031 1432
rect 3131 2208 3189 2220
rect 3131 1432 3143 2208
rect 3177 1432 3189 2208
rect 3131 1420 3189 1432
rect 3289 2208 3347 2220
rect 3289 1432 3301 2208
rect 3335 1432 3347 2208
rect 3289 1420 3347 1432
rect 3447 2208 3505 2220
rect 3447 1432 3459 2208
rect 3493 1432 3505 2208
rect 3447 1420 3505 1432
rect 3605 2208 3663 2220
rect 3605 1432 3617 2208
rect 3651 1432 3663 2208
rect 3605 1420 3663 1432
rect 3763 2208 3821 2220
rect 3763 1432 3775 2208
rect 3809 1432 3821 2208
rect 3763 1420 3821 1432
rect 3921 2208 3979 2220
rect 3921 1432 3933 2208
rect 3967 1432 3979 2208
rect 3921 1420 3979 1432
rect 4079 2208 4137 2220
rect 4079 1432 4091 2208
rect 4125 1432 4137 2208
rect 4079 1420 4137 1432
rect 4237 2208 4295 2220
rect 4237 1432 4249 2208
rect 4283 1432 4295 2208
rect 4237 1420 4295 1432
rect 4395 2208 4453 2220
rect 4395 1432 4407 2208
rect 4441 1432 4453 2208
rect 4395 1420 4453 1432
rect 4553 2208 4611 2220
rect 4553 1432 4565 2208
rect 4599 1432 4611 2208
rect 4553 1420 4611 1432
rect 4711 2208 4769 2220
rect 4711 1432 4723 2208
rect 4757 1432 4769 2208
rect 4711 1420 4769 1432
rect 4869 2208 4927 2220
rect 4869 1432 4881 2208
rect 4915 1432 4927 2208
rect 4869 1420 4927 1432
rect 5027 2208 5085 2220
rect 5027 1432 5039 2208
rect 5073 1432 5085 2208
rect 5027 1420 5085 1432
rect 5185 2208 5243 2220
rect 5185 1432 5197 2208
rect 5231 1432 5243 2208
rect 5185 1420 5243 1432
rect 5343 2208 5401 2220
rect 5343 1432 5355 2208
rect 5389 1432 5401 2208
rect 5343 1420 5401 1432
rect 5501 2208 5559 2220
rect 5501 1432 5513 2208
rect 5547 1432 5559 2208
rect 5501 1420 5559 1432
rect 5659 2208 5717 2220
rect 5659 1432 5671 2208
rect 5705 1432 5717 2208
rect 5659 1420 5717 1432
rect 5817 2208 5875 2220
rect 5817 1432 5829 2208
rect 5863 1432 5875 2208
rect 5817 1420 5875 1432
rect 5975 2208 6033 2220
rect 5975 1432 5987 2208
rect 6021 1432 6033 2208
rect 5975 1420 6033 1432
rect 6133 2208 6191 2220
rect 6133 1432 6145 2208
rect 6179 1432 6191 2208
rect 6133 1420 6191 1432
rect 6291 2208 6349 2220
rect 6291 1432 6303 2208
rect 6337 1432 6349 2208
rect 6291 1420 6349 1432
rect -6349 1298 -6291 1310
rect -6349 522 -6337 1298
rect -6303 522 -6291 1298
rect -6349 510 -6291 522
rect -6191 1298 -6133 1310
rect -6191 522 -6179 1298
rect -6145 522 -6133 1298
rect -6191 510 -6133 522
rect -6033 1298 -5975 1310
rect -6033 522 -6021 1298
rect -5987 522 -5975 1298
rect -6033 510 -5975 522
rect -5875 1298 -5817 1310
rect -5875 522 -5863 1298
rect -5829 522 -5817 1298
rect -5875 510 -5817 522
rect -5717 1298 -5659 1310
rect -5717 522 -5705 1298
rect -5671 522 -5659 1298
rect -5717 510 -5659 522
rect -5559 1298 -5501 1310
rect -5559 522 -5547 1298
rect -5513 522 -5501 1298
rect -5559 510 -5501 522
rect -5401 1298 -5343 1310
rect -5401 522 -5389 1298
rect -5355 522 -5343 1298
rect -5401 510 -5343 522
rect -5243 1298 -5185 1310
rect -5243 522 -5231 1298
rect -5197 522 -5185 1298
rect -5243 510 -5185 522
rect -5085 1298 -5027 1310
rect -5085 522 -5073 1298
rect -5039 522 -5027 1298
rect -5085 510 -5027 522
rect -4927 1298 -4869 1310
rect -4927 522 -4915 1298
rect -4881 522 -4869 1298
rect -4927 510 -4869 522
rect -4769 1298 -4711 1310
rect -4769 522 -4757 1298
rect -4723 522 -4711 1298
rect -4769 510 -4711 522
rect -4611 1298 -4553 1310
rect -4611 522 -4599 1298
rect -4565 522 -4553 1298
rect -4611 510 -4553 522
rect -4453 1298 -4395 1310
rect -4453 522 -4441 1298
rect -4407 522 -4395 1298
rect -4453 510 -4395 522
rect -4295 1298 -4237 1310
rect -4295 522 -4283 1298
rect -4249 522 -4237 1298
rect -4295 510 -4237 522
rect -4137 1298 -4079 1310
rect -4137 522 -4125 1298
rect -4091 522 -4079 1298
rect -4137 510 -4079 522
rect -3979 1298 -3921 1310
rect -3979 522 -3967 1298
rect -3933 522 -3921 1298
rect -3979 510 -3921 522
rect -3821 1298 -3763 1310
rect -3821 522 -3809 1298
rect -3775 522 -3763 1298
rect -3821 510 -3763 522
rect -3663 1298 -3605 1310
rect -3663 522 -3651 1298
rect -3617 522 -3605 1298
rect -3663 510 -3605 522
rect -3505 1298 -3447 1310
rect -3505 522 -3493 1298
rect -3459 522 -3447 1298
rect -3505 510 -3447 522
rect -3347 1298 -3289 1310
rect -3347 522 -3335 1298
rect -3301 522 -3289 1298
rect -3347 510 -3289 522
rect -3189 1298 -3131 1310
rect -3189 522 -3177 1298
rect -3143 522 -3131 1298
rect -3189 510 -3131 522
rect -3031 1298 -2973 1310
rect -3031 522 -3019 1298
rect -2985 522 -2973 1298
rect -3031 510 -2973 522
rect -2873 1298 -2815 1310
rect -2873 522 -2861 1298
rect -2827 522 -2815 1298
rect -2873 510 -2815 522
rect -2715 1298 -2657 1310
rect -2715 522 -2703 1298
rect -2669 522 -2657 1298
rect -2715 510 -2657 522
rect -2557 1298 -2499 1310
rect -2557 522 -2545 1298
rect -2511 522 -2499 1298
rect -2557 510 -2499 522
rect -2399 1298 -2341 1310
rect -2399 522 -2387 1298
rect -2353 522 -2341 1298
rect -2399 510 -2341 522
rect -2241 1298 -2183 1310
rect -2241 522 -2229 1298
rect -2195 522 -2183 1298
rect -2241 510 -2183 522
rect -2083 1298 -2025 1310
rect -2083 522 -2071 1298
rect -2037 522 -2025 1298
rect -2083 510 -2025 522
rect -1925 1298 -1867 1310
rect -1925 522 -1913 1298
rect -1879 522 -1867 1298
rect -1925 510 -1867 522
rect -1767 1298 -1709 1310
rect -1767 522 -1755 1298
rect -1721 522 -1709 1298
rect -1767 510 -1709 522
rect -1609 1298 -1551 1310
rect -1609 522 -1597 1298
rect -1563 522 -1551 1298
rect -1609 510 -1551 522
rect -1451 1298 -1393 1310
rect -1451 522 -1439 1298
rect -1405 522 -1393 1298
rect -1451 510 -1393 522
rect -1293 1298 -1235 1310
rect -1293 522 -1281 1298
rect -1247 522 -1235 1298
rect -1293 510 -1235 522
rect -1135 1298 -1077 1310
rect -1135 522 -1123 1298
rect -1089 522 -1077 1298
rect -1135 510 -1077 522
rect -977 1298 -919 1310
rect -977 522 -965 1298
rect -931 522 -919 1298
rect -977 510 -919 522
rect -819 1298 -761 1310
rect -819 522 -807 1298
rect -773 522 -761 1298
rect -819 510 -761 522
rect -661 1298 -603 1310
rect -661 522 -649 1298
rect -615 522 -603 1298
rect -661 510 -603 522
rect -503 1298 -445 1310
rect -503 522 -491 1298
rect -457 522 -445 1298
rect -503 510 -445 522
rect -345 1298 -287 1310
rect -345 522 -333 1298
rect -299 522 -287 1298
rect -345 510 -287 522
rect -187 1298 -129 1310
rect -187 522 -175 1298
rect -141 522 -129 1298
rect -187 510 -129 522
rect -29 1298 29 1310
rect -29 522 -17 1298
rect 17 522 29 1298
rect -29 510 29 522
rect 129 1298 187 1310
rect 129 522 141 1298
rect 175 522 187 1298
rect 129 510 187 522
rect 287 1298 345 1310
rect 287 522 299 1298
rect 333 522 345 1298
rect 287 510 345 522
rect 445 1298 503 1310
rect 445 522 457 1298
rect 491 522 503 1298
rect 445 510 503 522
rect 603 1298 661 1310
rect 603 522 615 1298
rect 649 522 661 1298
rect 603 510 661 522
rect 761 1298 819 1310
rect 761 522 773 1298
rect 807 522 819 1298
rect 761 510 819 522
rect 919 1298 977 1310
rect 919 522 931 1298
rect 965 522 977 1298
rect 919 510 977 522
rect 1077 1298 1135 1310
rect 1077 522 1089 1298
rect 1123 522 1135 1298
rect 1077 510 1135 522
rect 1235 1298 1293 1310
rect 1235 522 1247 1298
rect 1281 522 1293 1298
rect 1235 510 1293 522
rect 1393 1298 1451 1310
rect 1393 522 1405 1298
rect 1439 522 1451 1298
rect 1393 510 1451 522
rect 1551 1298 1609 1310
rect 1551 522 1563 1298
rect 1597 522 1609 1298
rect 1551 510 1609 522
rect 1709 1298 1767 1310
rect 1709 522 1721 1298
rect 1755 522 1767 1298
rect 1709 510 1767 522
rect 1867 1298 1925 1310
rect 1867 522 1879 1298
rect 1913 522 1925 1298
rect 1867 510 1925 522
rect 2025 1298 2083 1310
rect 2025 522 2037 1298
rect 2071 522 2083 1298
rect 2025 510 2083 522
rect 2183 1298 2241 1310
rect 2183 522 2195 1298
rect 2229 522 2241 1298
rect 2183 510 2241 522
rect 2341 1298 2399 1310
rect 2341 522 2353 1298
rect 2387 522 2399 1298
rect 2341 510 2399 522
rect 2499 1298 2557 1310
rect 2499 522 2511 1298
rect 2545 522 2557 1298
rect 2499 510 2557 522
rect 2657 1298 2715 1310
rect 2657 522 2669 1298
rect 2703 522 2715 1298
rect 2657 510 2715 522
rect 2815 1298 2873 1310
rect 2815 522 2827 1298
rect 2861 522 2873 1298
rect 2815 510 2873 522
rect 2973 1298 3031 1310
rect 2973 522 2985 1298
rect 3019 522 3031 1298
rect 2973 510 3031 522
rect 3131 1298 3189 1310
rect 3131 522 3143 1298
rect 3177 522 3189 1298
rect 3131 510 3189 522
rect 3289 1298 3347 1310
rect 3289 522 3301 1298
rect 3335 522 3347 1298
rect 3289 510 3347 522
rect 3447 1298 3505 1310
rect 3447 522 3459 1298
rect 3493 522 3505 1298
rect 3447 510 3505 522
rect 3605 1298 3663 1310
rect 3605 522 3617 1298
rect 3651 522 3663 1298
rect 3605 510 3663 522
rect 3763 1298 3821 1310
rect 3763 522 3775 1298
rect 3809 522 3821 1298
rect 3763 510 3821 522
rect 3921 1298 3979 1310
rect 3921 522 3933 1298
rect 3967 522 3979 1298
rect 3921 510 3979 522
rect 4079 1298 4137 1310
rect 4079 522 4091 1298
rect 4125 522 4137 1298
rect 4079 510 4137 522
rect 4237 1298 4295 1310
rect 4237 522 4249 1298
rect 4283 522 4295 1298
rect 4237 510 4295 522
rect 4395 1298 4453 1310
rect 4395 522 4407 1298
rect 4441 522 4453 1298
rect 4395 510 4453 522
rect 4553 1298 4611 1310
rect 4553 522 4565 1298
rect 4599 522 4611 1298
rect 4553 510 4611 522
rect 4711 1298 4769 1310
rect 4711 522 4723 1298
rect 4757 522 4769 1298
rect 4711 510 4769 522
rect 4869 1298 4927 1310
rect 4869 522 4881 1298
rect 4915 522 4927 1298
rect 4869 510 4927 522
rect 5027 1298 5085 1310
rect 5027 522 5039 1298
rect 5073 522 5085 1298
rect 5027 510 5085 522
rect 5185 1298 5243 1310
rect 5185 522 5197 1298
rect 5231 522 5243 1298
rect 5185 510 5243 522
rect 5343 1298 5401 1310
rect 5343 522 5355 1298
rect 5389 522 5401 1298
rect 5343 510 5401 522
rect 5501 1298 5559 1310
rect 5501 522 5513 1298
rect 5547 522 5559 1298
rect 5501 510 5559 522
rect 5659 1298 5717 1310
rect 5659 522 5671 1298
rect 5705 522 5717 1298
rect 5659 510 5717 522
rect 5817 1298 5875 1310
rect 5817 522 5829 1298
rect 5863 522 5875 1298
rect 5817 510 5875 522
rect 5975 1298 6033 1310
rect 5975 522 5987 1298
rect 6021 522 6033 1298
rect 5975 510 6033 522
rect 6133 1298 6191 1310
rect 6133 522 6145 1298
rect 6179 522 6191 1298
rect 6133 510 6191 522
rect 6291 1298 6349 1310
rect 6291 522 6303 1298
rect 6337 522 6349 1298
rect 6291 510 6349 522
rect -6349 388 -6291 400
rect -6349 -388 -6337 388
rect -6303 -388 -6291 388
rect -6349 -400 -6291 -388
rect -6191 388 -6133 400
rect -6191 -388 -6179 388
rect -6145 -388 -6133 388
rect -6191 -400 -6133 -388
rect -6033 388 -5975 400
rect -6033 -388 -6021 388
rect -5987 -388 -5975 388
rect -6033 -400 -5975 -388
rect -5875 388 -5817 400
rect -5875 -388 -5863 388
rect -5829 -388 -5817 388
rect -5875 -400 -5817 -388
rect -5717 388 -5659 400
rect -5717 -388 -5705 388
rect -5671 -388 -5659 388
rect -5717 -400 -5659 -388
rect -5559 388 -5501 400
rect -5559 -388 -5547 388
rect -5513 -388 -5501 388
rect -5559 -400 -5501 -388
rect -5401 388 -5343 400
rect -5401 -388 -5389 388
rect -5355 -388 -5343 388
rect -5401 -400 -5343 -388
rect -5243 388 -5185 400
rect -5243 -388 -5231 388
rect -5197 -388 -5185 388
rect -5243 -400 -5185 -388
rect -5085 388 -5027 400
rect -5085 -388 -5073 388
rect -5039 -388 -5027 388
rect -5085 -400 -5027 -388
rect -4927 388 -4869 400
rect -4927 -388 -4915 388
rect -4881 -388 -4869 388
rect -4927 -400 -4869 -388
rect -4769 388 -4711 400
rect -4769 -388 -4757 388
rect -4723 -388 -4711 388
rect -4769 -400 -4711 -388
rect -4611 388 -4553 400
rect -4611 -388 -4599 388
rect -4565 -388 -4553 388
rect -4611 -400 -4553 -388
rect -4453 388 -4395 400
rect -4453 -388 -4441 388
rect -4407 -388 -4395 388
rect -4453 -400 -4395 -388
rect -4295 388 -4237 400
rect -4295 -388 -4283 388
rect -4249 -388 -4237 388
rect -4295 -400 -4237 -388
rect -4137 388 -4079 400
rect -4137 -388 -4125 388
rect -4091 -388 -4079 388
rect -4137 -400 -4079 -388
rect -3979 388 -3921 400
rect -3979 -388 -3967 388
rect -3933 -388 -3921 388
rect -3979 -400 -3921 -388
rect -3821 388 -3763 400
rect -3821 -388 -3809 388
rect -3775 -388 -3763 388
rect -3821 -400 -3763 -388
rect -3663 388 -3605 400
rect -3663 -388 -3651 388
rect -3617 -388 -3605 388
rect -3663 -400 -3605 -388
rect -3505 388 -3447 400
rect -3505 -388 -3493 388
rect -3459 -388 -3447 388
rect -3505 -400 -3447 -388
rect -3347 388 -3289 400
rect -3347 -388 -3335 388
rect -3301 -388 -3289 388
rect -3347 -400 -3289 -388
rect -3189 388 -3131 400
rect -3189 -388 -3177 388
rect -3143 -388 -3131 388
rect -3189 -400 -3131 -388
rect -3031 388 -2973 400
rect -3031 -388 -3019 388
rect -2985 -388 -2973 388
rect -3031 -400 -2973 -388
rect -2873 388 -2815 400
rect -2873 -388 -2861 388
rect -2827 -388 -2815 388
rect -2873 -400 -2815 -388
rect -2715 388 -2657 400
rect -2715 -388 -2703 388
rect -2669 -388 -2657 388
rect -2715 -400 -2657 -388
rect -2557 388 -2499 400
rect -2557 -388 -2545 388
rect -2511 -388 -2499 388
rect -2557 -400 -2499 -388
rect -2399 388 -2341 400
rect -2399 -388 -2387 388
rect -2353 -388 -2341 388
rect -2399 -400 -2341 -388
rect -2241 388 -2183 400
rect -2241 -388 -2229 388
rect -2195 -388 -2183 388
rect -2241 -400 -2183 -388
rect -2083 388 -2025 400
rect -2083 -388 -2071 388
rect -2037 -388 -2025 388
rect -2083 -400 -2025 -388
rect -1925 388 -1867 400
rect -1925 -388 -1913 388
rect -1879 -388 -1867 388
rect -1925 -400 -1867 -388
rect -1767 388 -1709 400
rect -1767 -388 -1755 388
rect -1721 -388 -1709 388
rect -1767 -400 -1709 -388
rect -1609 388 -1551 400
rect -1609 -388 -1597 388
rect -1563 -388 -1551 388
rect -1609 -400 -1551 -388
rect -1451 388 -1393 400
rect -1451 -388 -1439 388
rect -1405 -388 -1393 388
rect -1451 -400 -1393 -388
rect -1293 388 -1235 400
rect -1293 -388 -1281 388
rect -1247 -388 -1235 388
rect -1293 -400 -1235 -388
rect -1135 388 -1077 400
rect -1135 -388 -1123 388
rect -1089 -388 -1077 388
rect -1135 -400 -1077 -388
rect -977 388 -919 400
rect -977 -388 -965 388
rect -931 -388 -919 388
rect -977 -400 -919 -388
rect -819 388 -761 400
rect -819 -388 -807 388
rect -773 -388 -761 388
rect -819 -400 -761 -388
rect -661 388 -603 400
rect -661 -388 -649 388
rect -615 -388 -603 388
rect -661 -400 -603 -388
rect -503 388 -445 400
rect -503 -388 -491 388
rect -457 -388 -445 388
rect -503 -400 -445 -388
rect -345 388 -287 400
rect -345 -388 -333 388
rect -299 -388 -287 388
rect -345 -400 -287 -388
rect -187 388 -129 400
rect -187 -388 -175 388
rect -141 -388 -129 388
rect -187 -400 -129 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 129 388 187 400
rect 129 -388 141 388
rect 175 -388 187 388
rect 129 -400 187 -388
rect 287 388 345 400
rect 287 -388 299 388
rect 333 -388 345 388
rect 287 -400 345 -388
rect 445 388 503 400
rect 445 -388 457 388
rect 491 -388 503 388
rect 445 -400 503 -388
rect 603 388 661 400
rect 603 -388 615 388
rect 649 -388 661 388
rect 603 -400 661 -388
rect 761 388 819 400
rect 761 -388 773 388
rect 807 -388 819 388
rect 761 -400 819 -388
rect 919 388 977 400
rect 919 -388 931 388
rect 965 -388 977 388
rect 919 -400 977 -388
rect 1077 388 1135 400
rect 1077 -388 1089 388
rect 1123 -388 1135 388
rect 1077 -400 1135 -388
rect 1235 388 1293 400
rect 1235 -388 1247 388
rect 1281 -388 1293 388
rect 1235 -400 1293 -388
rect 1393 388 1451 400
rect 1393 -388 1405 388
rect 1439 -388 1451 388
rect 1393 -400 1451 -388
rect 1551 388 1609 400
rect 1551 -388 1563 388
rect 1597 -388 1609 388
rect 1551 -400 1609 -388
rect 1709 388 1767 400
rect 1709 -388 1721 388
rect 1755 -388 1767 388
rect 1709 -400 1767 -388
rect 1867 388 1925 400
rect 1867 -388 1879 388
rect 1913 -388 1925 388
rect 1867 -400 1925 -388
rect 2025 388 2083 400
rect 2025 -388 2037 388
rect 2071 -388 2083 388
rect 2025 -400 2083 -388
rect 2183 388 2241 400
rect 2183 -388 2195 388
rect 2229 -388 2241 388
rect 2183 -400 2241 -388
rect 2341 388 2399 400
rect 2341 -388 2353 388
rect 2387 -388 2399 388
rect 2341 -400 2399 -388
rect 2499 388 2557 400
rect 2499 -388 2511 388
rect 2545 -388 2557 388
rect 2499 -400 2557 -388
rect 2657 388 2715 400
rect 2657 -388 2669 388
rect 2703 -388 2715 388
rect 2657 -400 2715 -388
rect 2815 388 2873 400
rect 2815 -388 2827 388
rect 2861 -388 2873 388
rect 2815 -400 2873 -388
rect 2973 388 3031 400
rect 2973 -388 2985 388
rect 3019 -388 3031 388
rect 2973 -400 3031 -388
rect 3131 388 3189 400
rect 3131 -388 3143 388
rect 3177 -388 3189 388
rect 3131 -400 3189 -388
rect 3289 388 3347 400
rect 3289 -388 3301 388
rect 3335 -388 3347 388
rect 3289 -400 3347 -388
rect 3447 388 3505 400
rect 3447 -388 3459 388
rect 3493 -388 3505 388
rect 3447 -400 3505 -388
rect 3605 388 3663 400
rect 3605 -388 3617 388
rect 3651 -388 3663 388
rect 3605 -400 3663 -388
rect 3763 388 3821 400
rect 3763 -388 3775 388
rect 3809 -388 3821 388
rect 3763 -400 3821 -388
rect 3921 388 3979 400
rect 3921 -388 3933 388
rect 3967 -388 3979 388
rect 3921 -400 3979 -388
rect 4079 388 4137 400
rect 4079 -388 4091 388
rect 4125 -388 4137 388
rect 4079 -400 4137 -388
rect 4237 388 4295 400
rect 4237 -388 4249 388
rect 4283 -388 4295 388
rect 4237 -400 4295 -388
rect 4395 388 4453 400
rect 4395 -388 4407 388
rect 4441 -388 4453 388
rect 4395 -400 4453 -388
rect 4553 388 4611 400
rect 4553 -388 4565 388
rect 4599 -388 4611 388
rect 4553 -400 4611 -388
rect 4711 388 4769 400
rect 4711 -388 4723 388
rect 4757 -388 4769 388
rect 4711 -400 4769 -388
rect 4869 388 4927 400
rect 4869 -388 4881 388
rect 4915 -388 4927 388
rect 4869 -400 4927 -388
rect 5027 388 5085 400
rect 5027 -388 5039 388
rect 5073 -388 5085 388
rect 5027 -400 5085 -388
rect 5185 388 5243 400
rect 5185 -388 5197 388
rect 5231 -388 5243 388
rect 5185 -400 5243 -388
rect 5343 388 5401 400
rect 5343 -388 5355 388
rect 5389 -388 5401 388
rect 5343 -400 5401 -388
rect 5501 388 5559 400
rect 5501 -388 5513 388
rect 5547 -388 5559 388
rect 5501 -400 5559 -388
rect 5659 388 5717 400
rect 5659 -388 5671 388
rect 5705 -388 5717 388
rect 5659 -400 5717 -388
rect 5817 388 5875 400
rect 5817 -388 5829 388
rect 5863 -388 5875 388
rect 5817 -400 5875 -388
rect 5975 388 6033 400
rect 5975 -388 5987 388
rect 6021 -388 6033 388
rect 5975 -400 6033 -388
rect 6133 388 6191 400
rect 6133 -388 6145 388
rect 6179 -388 6191 388
rect 6133 -400 6191 -388
rect 6291 388 6349 400
rect 6291 -388 6303 388
rect 6337 -388 6349 388
rect 6291 -400 6349 -388
rect -6349 -522 -6291 -510
rect -6349 -1298 -6337 -522
rect -6303 -1298 -6291 -522
rect -6349 -1310 -6291 -1298
rect -6191 -522 -6133 -510
rect -6191 -1298 -6179 -522
rect -6145 -1298 -6133 -522
rect -6191 -1310 -6133 -1298
rect -6033 -522 -5975 -510
rect -6033 -1298 -6021 -522
rect -5987 -1298 -5975 -522
rect -6033 -1310 -5975 -1298
rect -5875 -522 -5817 -510
rect -5875 -1298 -5863 -522
rect -5829 -1298 -5817 -522
rect -5875 -1310 -5817 -1298
rect -5717 -522 -5659 -510
rect -5717 -1298 -5705 -522
rect -5671 -1298 -5659 -522
rect -5717 -1310 -5659 -1298
rect -5559 -522 -5501 -510
rect -5559 -1298 -5547 -522
rect -5513 -1298 -5501 -522
rect -5559 -1310 -5501 -1298
rect -5401 -522 -5343 -510
rect -5401 -1298 -5389 -522
rect -5355 -1298 -5343 -522
rect -5401 -1310 -5343 -1298
rect -5243 -522 -5185 -510
rect -5243 -1298 -5231 -522
rect -5197 -1298 -5185 -522
rect -5243 -1310 -5185 -1298
rect -5085 -522 -5027 -510
rect -5085 -1298 -5073 -522
rect -5039 -1298 -5027 -522
rect -5085 -1310 -5027 -1298
rect -4927 -522 -4869 -510
rect -4927 -1298 -4915 -522
rect -4881 -1298 -4869 -522
rect -4927 -1310 -4869 -1298
rect -4769 -522 -4711 -510
rect -4769 -1298 -4757 -522
rect -4723 -1298 -4711 -522
rect -4769 -1310 -4711 -1298
rect -4611 -522 -4553 -510
rect -4611 -1298 -4599 -522
rect -4565 -1298 -4553 -522
rect -4611 -1310 -4553 -1298
rect -4453 -522 -4395 -510
rect -4453 -1298 -4441 -522
rect -4407 -1298 -4395 -522
rect -4453 -1310 -4395 -1298
rect -4295 -522 -4237 -510
rect -4295 -1298 -4283 -522
rect -4249 -1298 -4237 -522
rect -4295 -1310 -4237 -1298
rect -4137 -522 -4079 -510
rect -4137 -1298 -4125 -522
rect -4091 -1298 -4079 -522
rect -4137 -1310 -4079 -1298
rect -3979 -522 -3921 -510
rect -3979 -1298 -3967 -522
rect -3933 -1298 -3921 -522
rect -3979 -1310 -3921 -1298
rect -3821 -522 -3763 -510
rect -3821 -1298 -3809 -522
rect -3775 -1298 -3763 -522
rect -3821 -1310 -3763 -1298
rect -3663 -522 -3605 -510
rect -3663 -1298 -3651 -522
rect -3617 -1298 -3605 -522
rect -3663 -1310 -3605 -1298
rect -3505 -522 -3447 -510
rect -3505 -1298 -3493 -522
rect -3459 -1298 -3447 -522
rect -3505 -1310 -3447 -1298
rect -3347 -522 -3289 -510
rect -3347 -1298 -3335 -522
rect -3301 -1298 -3289 -522
rect -3347 -1310 -3289 -1298
rect -3189 -522 -3131 -510
rect -3189 -1298 -3177 -522
rect -3143 -1298 -3131 -522
rect -3189 -1310 -3131 -1298
rect -3031 -522 -2973 -510
rect -3031 -1298 -3019 -522
rect -2985 -1298 -2973 -522
rect -3031 -1310 -2973 -1298
rect -2873 -522 -2815 -510
rect -2873 -1298 -2861 -522
rect -2827 -1298 -2815 -522
rect -2873 -1310 -2815 -1298
rect -2715 -522 -2657 -510
rect -2715 -1298 -2703 -522
rect -2669 -1298 -2657 -522
rect -2715 -1310 -2657 -1298
rect -2557 -522 -2499 -510
rect -2557 -1298 -2545 -522
rect -2511 -1298 -2499 -522
rect -2557 -1310 -2499 -1298
rect -2399 -522 -2341 -510
rect -2399 -1298 -2387 -522
rect -2353 -1298 -2341 -522
rect -2399 -1310 -2341 -1298
rect -2241 -522 -2183 -510
rect -2241 -1298 -2229 -522
rect -2195 -1298 -2183 -522
rect -2241 -1310 -2183 -1298
rect -2083 -522 -2025 -510
rect -2083 -1298 -2071 -522
rect -2037 -1298 -2025 -522
rect -2083 -1310 -2025 -1298
rect -1925 -522 -1867 -510
rect -1925 -1298 -1913 -522
rect -1879 -1298 -1867 -522
rect -1925 -1310 -1867 -1298
rect -1767 -522 -1709 -510
rect -1767 -1298 -1755 -522
rect -1721 -1298 -1709 -522
rect -1767 -1310 -1709 -1298
rect -1609 -522 -1551 -510
rect -1609 -1298 -1597 -522
rect -1563 -1298 -1551 -522
rect -1609 -1310 -1551 -1298
rect -1451 -522 -1393 -510
rect -1451 -1298 -1439 -522
rect -1405 -1298 -1393 -522
rect -1451 -1310 -1393 -1298
rect -1293 -522 -1235 -510
rect -1293 -1298 -1281 -522
rect -1247 -1298 -1235 -522
rect -1293 -1310 -1235 -1298
rect -1135 -522 -1077 -510
rect -1135 -1298 -1123 -522
rect -1089 -1298 -1077 -522
rect -1135 -1310 -1077 -1298
rect -977 -522 -919 -510
rect -977 -1298 -965 -522
rect -931 -1298 -919 -522
rect -977 -1310 -919 -1298
rect -819 -522 -761 -510
rect -819 -1298 -807 -522
rect -773 -1298 -761 -522
rect -819 -1310 -761 -1298
rect -661 -522 -603 -510
rect -661 -1298 -649 -522
rect -615 -1298 -603 -522
rect -661 -1310 -603 -1298
rect -503 -522 -445 -510
rect -503 -1298 -491 -522
rect -457 -1298 -445 -522
rect -503 -1310 -445 -1298
rect -345 -522 -287 -510
rect -345 -1298 -333 -522
rect -299 -1298 -287 -522
rect -345 -1310 -287 -1298
rect -187 -522 -129 -510
rect -187 -1298 -175 -522
rect -141 -1298 -129 -522
rect -187 -1310 -129 -1298
rect -29 -522 29 -510
rect -29 -1298 -17 -522
rect 17 -1298 29 -522
rect -29 -1310 29 -1298
rect 129 -522 187 -510
rect 129 -1298 141 -522
rect 175 -1298 187 -522
rect 129 -1310 187 -1298
rect 287 -522 345 -510
rect 287 -1298 299 -522
rect 333 -1298 345 -522
rect 287 -1310 345 -1298
rect 445 -522 503 -510
rect 445 -1298 457 -522
rect 491 -1298 503 -522
rect 445 -1310 503 -1298
rect 603 -522 661 -510
rect 603 -1298 615 -522
rect 649 -1298 661 -522
rect 603 -1310 661 -1298
rect 761 -522 819 -510
rect 761 -1298 773 -522
rect 807 -1298 819 -522
rect 761 -1310 819 -1298
rect 919 -522 977 -510
rect 919 -1298 931 -522
rect 965 -1298 977 -522
rect 919 -1310 977 -1298
rect 1077 -522 1135 -510
rect 1077 -1298 1089 -522
rect 1123 -1298 1135 -522
rect 1077 -1310 1135 -1298
rect 1235 -522 1293 -510
rect 1235 -1298 1247 -522
rect 1281 -1298 1293 -522
rect 1235 -1310 1293 -1298
rect 1393 -522 1451 -510
rect 1393 -1298 1405 -522
rect 1439 -1298 1451 -522
rect 1393 -1310 1451 -1298
rect 1551 -522 1609 -510
rect 1551 -1298 1563 -522
rect 1597 -1298 1609 -522
rect 1551 -1310 1609 -1298
rect 1709 -522 1767 -510
rect 1709 -1298 1721 -522
rect 1755 -1298 1767 -522
rect 1709 -1310 1767 -1298
rect 1867 -522 1925 -510
rect 1867 -1298 1879 -522
rect 1913 -1298 1925 -522
rect 1867 -1310 1925 -1298
rect 2025 -522 2083 -510
rect 2025 -1298 2037 -522
rect 2071 -1298 2083 -522
rect 2025 -1310 2083 -1298
rect 2183 -522 2241 -510
rect 2183 -1298 2195 -522
rect 2229 -1298 2241 -522
rect 2183 -1310 2241 -1298
rect 2341 -522 2399 -510
rect 2341 -1298 2353 -522
rect 2387 -1298 2399 -522
rect 2341 -1310 2399 -1298
rect 2499 -522 2557 -510
rect 2499 -1298 2511 -522
rect 2545 -1298 2557 -522
rect 2499 -1310 2557 -1298
rect 2657 -522 2715 -510
rect 2657 -1298 2669 -522
rect 2703 -1298 2715 -522
rect 2657 -1310 2715 -1298
rect 2815 -522 2873 -510
rect 2815 -1298 2827 -522
rect 2861 -1298 2873 -522
rect 2815 -1310 2873 -1298
rect 2973 -522 3031 -510
rect 2973 -1298 2985 -522
rect 3019 -1298 3031 -522
rect 2973 -1310 3031 -1298
rect 3131 -522 3189 -510
rect 3131 -1298 3143 -522
rect 3177 -1298 3189 -522
rect 3131 -1310 3189 -1298
rect 3289 -522 3347 -510
rect 3289 -1298 3301 -522
rect 3335 -1298 3347 -522
rect 3289 -1310 3347 -1298
rect 3447 -522 3505 -510
rect 3447 -1298 3459 -522
rect 3493 -1298 3505 -522
rect 3447 -1310 3505 -1298
rect 3605 -522 3663 -510
rect 3605 -1298 3617 -522
rect 3651 -1298 3663 -522
rect 3605 -1310 3663 -1298
rect 3763 -522 3821 -510
rect 3763 -1298 3775 -522
rect 3809 -1298 3821 -522
rect 3763 -1310 3821 -1298
rect 3921 -522 3979 -510
rect 3921 -1298 3933 -522
rect 3967 -1298 3979 -522
rect 3921 -1310 3979 -1298
rect 4079 -522 4137 -510
rect 4079 -1298 4091 -522
rect 4125 -1298 4137 -522
rect 4079 -1310 4137 -1298
rect 4237 -522 4295 -510
rect 4237 -1298 4249 -522
rect 4283 -1298 4295 -522
rect 4237 -1310 4295 -1298
rect 4395 -522 4453 -510
rect 4395 -1298 4407 -522
rect 4441 -1298 4453 -522
rect 4395 -1310 4453 -1298
rect 4553 -522 4611 -510
rect 4553 -1298 4565 -522
rect 4599 -1298 4611 -522
rect 4553 -1310 4611 -1298
rect 4711 -522 4769 -510
rect 4711 -1298 4723 -522
rect 4757 -1298 4769 -522
rect 4711 -1310 4769 -1298
rect 4869 -522 4927 -510
rect 4869 -1298 4881 -522
rect 4915 -1298 4927 -522
rect 4869 -1310 4927 -1298
rect 5027 -522 5085 -510
rect 5027 -1298 5039 -522
rect 5073 -1298 5085 -522
rect 5027 -1310 5085 -1298
rect 5185 -522 5243 -510
rect 5185 -1298 5197 -522
rect 5231 -1298 5243 -522
rect 5185 -1310 5243 -1298
rect 5343 -522 5401 -510
rect 5343 -1298 5355 -522
rect 5389 -1298 5401 -522
rect 5343 -1310 5401 -1298
rect 5501 -522 5559 -510
rect 5501 -1298 5513 -522
rect 5547 -1298 5559 -522
rect 5501 -1310 5559 -1298
rect 5659 -522 5717 -510
rect 5659 -1298 5671 -522
rect 5705 -1298 5717 -522
rect 5659 -1310 5717 -1298
rect 5817 -522 5875 -510
rect 5817 -1298 5829 -522
rect 5863 -1298 5875 -522
rect 5817 -1310 5875 -1298
rect 5975 -522 6033 -510
rect 5975 -1298 5987 -522
rect 6021 -1298 6033 -522
rect 5975 -1310 6033 -1298
rect 6133 -522 6191 -510
rect 6133 -1298 6145 -522
rect 6179 -1298 6191 -522
rect 6133 -1310 6191 -1298
rect 6291 -522 6349 -510
rect 6291 -1298 6303 -522
rect 6337 -1298 6349 -522
rect 6291 -1310 6349 -1298
rect -6349 -1432 -6291 -1420
rect -6349 -2208 -6337 -1432
rect -6303 -2208 -6291 -1432
rect -6349 -2220 -6291 -2208
rect -6191 -1432 -6133 -1420
rect -6191 -2208 -6179 -1432
rect -6145 -2208 -6133 -1432
rect -6191 -2220 -6133 -2208
rect -6033 -1432 -5975 -1420
rect -6033 -2208 -6021 -1432
rect -5987 -2208 -5975 -1432
rect -6033 -2220 -5975 -2208
rect -5875 -1432 -5817 -1420
rect -5875 -2208 -5863 -1432
rect -5829 -2208 -5817 -1432
rect -5875 -2220 -5817 -2208
rect -5717 -1432 -5659 -1420
rect -5717 -2208 -5705 -1432
rect -5671 -2208 -5659 -1432
rect -5717 -2220 -5659 -2208
rect -5559 -1432 -5501 -1420
rect -5559 -2208 -5547 -1432
rect -5513 -2208 -5501 -1432
rect -5559 -2220 -5501 -2208
rect -5401 -1432 -5343 -1420
rect -5401 -2208 -5389 -1432
rect -5355 -2208 -5343 -1432
rect -5401 -2220 -5343 -2208
rect -5243 -1432 -5185 -1420
rect -5243 -2208 -5231 -1432
rect -5197 -2208 -5185 -1432
rect -5243 -2220 -5185 -2208
rect -5085 -1432 -5027 -1420
rect -5085 -2208 -5073 -1432
rect -5039 -2208 -5027 -1432
rect -5085 -2220 -5027 -2208
rect -4927 -1432 -4869 -1420
rect -4927 -2208 -4915 -1432
rect -4881 -2208 -4869 -1432
rect -4927 -2220 -4869 -2208
rect -4769 -1432 -4711 -1420
rect -4769 -2208 -4757 -1432
rect -4723 -2208 -4711 -1432
rect -4769 -2220 -4711 -2208
rect -4611 -1432 -4553 -1420
rect -4611 -2208 -4599 -1432
rect -4565 -2208 -4553 -1432
rect -4611 -2220 -4553 -2208
rect -4453 -1432 -4395 -1420
rect -4453 -2208 -4441 -1432
rect -4407 -2208 -4395 -1432
rect -4453 -2220 -4395 -2208
rect -4295 -1432 -4237 -1420
rect -4295 -2208 -4283 -1432
rect -4249 -2208 -4237 -1432
rect -4295 -2220 -4237 -2208
rect -4137 -1432 -4079 -1420
rect -4137 -2208 -4125 -1432
rect -4091 -2208 -4079 -1432
rect -4137 -2220 -4079 -2208
rect -3979 -1432 -3921 -1420
rect -3979 -2208 -3967 -1432
rect -3933 -2208 -3921 -1432
rect -3979 -2220 -3921 -2208
rect -3821 -1432 -3763 -1420
rect -3821 -2208 -3809 -1432
rect -3775 -2208 -3763 -1432
rect -3821 -2220 -3763 -2208
rect -3663 -1432 -3605 -1420
rect -3663 -2208 -3651 -1432
rect -3617 -2208 -3605 -1432
rect -3663 -2220 -3605 -2208
rect -3505 -1432 -3447 -1420
rect -3505 -2208 -3493 -1432
rect -3459 -2208 -3447 -1432
rect -3505 -2220 -3447 -2208
rect -3347 -1432 -3289 -1420
rect -3347 -2208 -3335 -1432
rect -3301 -2208 -3289 -1432
rect -3347 -2220 -3289 -2208
rect -3189 -1432 -3131 -1420
rect -3189 -2208 -3177 -1432
rect -3143 -2208 -3131 -1432
rect -3189 -2220 -3131 -2208
rect -3031 -1432 -2973 -1420
rect -3031 -2208 -3019 -1432
rect -2985 -2208 -2973 -1432
rect -3031 -2220 -2973 -2208
rect -2873 -1432 -2815 -1420
rect -2873 -2208 -2861 -1432
rect -2827 -2208 -2815 -1432
rect -2873 -2220 -2815 -2208
rect -2715 -1432 -2657 -1420
rect -2715 -2208 -2703 -1432
rect -2669 -2208 -2657 -1432
rect -2715 -2220 -2657 -2208
rect -2557 -1432 -2499 -1420
rect -2557 -2208 -2545 -1432
rect -2511 -2208 -2499 -1432
rect -2557 -2220 -2499 -2208
rect -2399 -1432 -2341 -1420
rect -2399 -2208 -2387 -1432
rect -2353 -2208 -2341 -1432
rect -2399 -2220 -2341 -2208
rect -2241 -1432 -2183 -1420
rect -2241 -2208 -2229 -1432
rect -2195 -2208 -2183 -1432
rect -2241 -2220 -2183 -2208
rect -2083 -1432 -2025 -1420
rect -2083 -2208 -2071 -1432
rect -2037 -2208 -2025 -1432
rect -2083 -2220 -2025 -2208
rect -1925 -1432 -1867 -1420
rect -1925 -2208 -1913 -1432
rect -1879 -2208 -1867 -1432
rect -1925 -2220 -1867 -2208
rect -1767 -1432 -1709 -1420
rect -1767 -2208 -1755 -1432
rect -1721 -2208 -1709 -1432
rect -1767 -2220 -1709 -2208
rect -1609 -1432 -1551 -1420
rect -1609 -2208 -1597 -1432
rect -1563 -2208 -1551 -1432
rect -1609 -2220 -1551 -2208
rect -1451 -1432 -1393 -1420
rect -1451 -2208 -1439 -1432
rect -1405 -2208 -1393 -1432
rect -1451 -2220 -1393 -2208
rect -1293 -1432 -1235 -1420
rect -1293 -2208 -1281 -1432
rect -1247 -2208 -1235 -1432
rect -1293 -2220 -1235 -2208
rect -1135 -1432 -1077 -1420
rect -1135 -2208 -1123 -1432
rect -1089 -2208 -1077 -1432
rect -1135 -2220 -1077 -2208
rect -977 -1432 -919 -1420
rect -977 -2208 -965 -1432
rect -931 -2208 -919 -1432
rect -977 -2220 -919 -2208
rect -819 -1432 -761 -1420
rect -819 -2208 -807 -1432
rect -773 -2208 -761 -1432
rect -819 -2220 -761 -2208
rect -661 -1432 -603 -1420
rect -661 -2208 -649 -1432
rect -615 -2208 -603 -1432
rect -661 -2220 -603 -2208
rect -503 -1432 -445 -1420
rect -503 -2208 -491 -1432
rect -457 -2208 -445 -1432
rect -503 -2220 -445 -2208
rect -345 -1432 -287 -1420
rect -345 -2208 -333 -1432
rect -299 -2208 -287 -1432
rect -345 -2220 -287 -2208
rect -187 -1432 -129 -1420
rect -187 -2208 -175 -1432
rect -141 -2208 -129 -1432
rect -187 -2220 -129 -2208
rect -29 -1432 29 -1420
rect -29 -2208 -17 -1432
rect 17 -2208 29 -1432
rect -29 -2220 29 -2208
rect 129 -1432 187 -1420
rect 129 -2208 141 -1432
rect 175 -2208 187 -1432
rect 129 -2220 187 -2208
rect 287 -1432 345 -1420
rect 287 -2208 299 -1432
rect 333 -2208 345 -1432
rect 287 -2220 345 -2208
rect 445 -1432 503 -1420
rect 445 -2208 457 -1432
rect 491 -2208 503 -1432
rect 445 -2220 503 -2208
rect 603 -1432 661 -1420
rect 603 -2208 615 -1432
rect 649 -2208 661 -1432
rect 603 -2220 661 -2208
rect 761 -1432 819 -1420
rect 761 -2208 773 -1432
rect 807 -2208 819 -1432
rect 761 -2220 819 -2208
rect 919 -1432 977 -1420
rect 919 -2208 931 -1432
rect 965 -2208 977 -1432
rect 919 -2220 977 -2208
rect 1077 -1432 1135 -1420
rect 1077 -2208 1089 -1432
rect 1123 -2208 1135 -1432
rect 1077 -2220 1135 -2208
rect 1235 -1432 1293 -1420
rect 1235 -2208 1247 -1432
rect 1281 -2208 1293 -1432
rect 1235 -2220 1293 -2208
rect 1393 -1432 1451 -1420
rect 1393 -2208 1405 -1432
rect 1439 -2208 1451 -1432
rect 1393 -2220 1451 -2208
rect 1551 -1432 1609 -1420
rect 1551 -2208 1563 -1432
rect 1597 -2208 1609 -1432
rect 1551 -2220 1609 -2208
rect 1709 -1432 1767 -1420
rect 1709 -2208 1721 -1432
rect 1755 -2208 1767 -1432
rect 1709 -2220 1767 -2208
rect 1867 -1432 1925 -1420
rect 1867 -2208 1879 -1432
rect 1913 -2208 1925 -1432
rect 1867 -2220 1925 -2208
rect 2025 -1432 2083 -1420
rect 2025 -2208 2037 -1432
rect 2071 -2208 2083 -1432
rect 2025 -2220 2083 -2208
rect 2183 -1432 2241 -1420
rect 2183 -2208 2195 -1432
rect 2229 -2208 2241 -1432
rect 2183 -2220 2241 -2208
rect 2341 -1432 2399 -1420
rect 2341 -2208 2353 -1432
rect 2387 -2208 2399 -1432
rect 2341 -2220 2399 -2208
rect 2499 -1432 2557 -1420
rect 2499 -2208 2511 -1432
rect 2545 -2208 2557 -1432
rect 2499 -2220 2557 -2208
rect 2657 -1432 2715 -1420
rect 2657 -2208 2669 -1432
rect 2703 -2208 2715 -1432
rect 2657 -2220 2715 -2208
rect 2815 -1432 2873 -1420
rect 2815 -2208 2827 -1432
rect 2861 -2208 2873 -1432
rect 2815 -2220 2873 -2208
rect 2973 -1432 3031 -1420
rect 2973 -2208 2985 -1432
rect 3019 -2208 3031 -1432
rect 2973 -2220 3031 -2208
rect 3131 -1432 3189 -1420
rect 3131 -2208 3143 -1432
rect 3177 -2208 3189 -1432
rect 3131 -2220 3189 -2208
rect 3289 -1432 3347 -1420
rect 3289 -2208 3301 -1432
rect 3335 -2208 3347 -1432
rect 3289 -2220 3347 -2208
rect 3447 -1432 3505 -1420
rect 3447 -2208 3459 -1432
rect 3493 -2208 3505 -1432
rect 3447 -2220 3505 -2208
rect 3605 -1432 3663 -1420
rect 3605 -2208 3617 -1432
rect 3651 -2208 3663 -1432
rect 3605 -2220 3663 -2208
rect 3763 -1432 3821 -1420
rect 3763 -2208 3775 -1432
rect 3809 -2208 3821 -1432
rect 3763 -2220 3821 -2208
rect 3921 -1432 3979 -1420
rect 3921 -2208 3933 -1432
rect 3967 -2208 3979 -1432
rect 3921 -2220 3979 -2208
rect 4079 -1432 4137 -1420
rect 4079 -2208 4091 -1432
rect 4125 -2208 4137 -1432
rect 4079 -2220 4137 -2208
rect 4237 -1432 4295 -1420
rect 4237 -2208 4249 -1432
rect 4283 -2208 4295 -1432
rect 4237 -2220 4295 -2208
rect 4395 -1432 4453 -1420
rect 4395 -2208 4407 -1432
rect 4441 -2208 4453 -1432
rect 4395 -2220 4453 -2208
rect 4553 -1432 4611 -1420
rect 4553 -2208 4565 -1432
rect 4599 -2208 4611 -1432
rect 4553 -2220 4611 -2208
rect 4711 -1432 4769 -1420
rect 4711 -2208 4723 -1432
rect 4757 -2208 4769 -1432
rect 4711 -2220 4769 -2208
rect 4869 -1432 4927 -1420
rect 4869 -2208 4881 -1432
rect 4915 -2208 4927 -1432
rect 4869 -2220 4927 -2208
rect 5027 -1432 5085 -1420
rect 5027 -2208 5039 -1432
rect 5073 -2208 5085 -1432
rect 5027 -2220 5085 -2208
rect 5185 -1432 5243 -1420
rect 5185 -2208 5197 -1432
rect 5231 -2208 5243 -1432
rect 5185 -2220 5243 -2208
rect 5343 -1432 5401 -1420
rect 5343 -2208 5355 -1432
rect 5389 -2208 5401 -1432
rect 5343 -2220 5401 -2208
rect 5501 -1432 5559 -1420
rect 5501 -2208 5513 -1432
rect 5547 -2208 5559 -1432
rect 5501 -2220 5559 -2208
rect 5659 -1432 5717 -1420
rect 5659 -2208 5671 -1432
rect 5705 -2208 5717 -1432
rect 5659 -2220 5717 -2208
rect 5817 -1432 5875 -1420
rect 5817 -2208 5829 -1432
rect 5863 -2208 5875 -1432
rect 5817 -2220 5875 -2208
rect 5975 -1432 6033 -1420
rect 5975 -2208 5987 -1432
rect 6021 -2208 6033 -1432
rect 5975 -2220 6033 -2208
rect 6133 -1432 6191 -1420
rect 6133 -2208 6145 -1432
rect 6179 -2208 6191 -1432
rect 6133 -2220 6191 -2208
rect 6291 -1432 6349 -1420
rect 6291 -2208 6303 -1432
rect 6337 -2208 6349 -1432
rect 6291 -2220 6349 -2208
<< mvndiffc >>
rect -6337 1432 -6303 2208
rect -6179 1432 -6145 2208
rect -6021 1432 -5987 2208
rect -5863 1432 -5829 2208
rect -5705 1432 -5671 2208
rect -5547 1432 -5513 2208
rect -5389 1432 -5355 2208
rect -5231 1432 -5197 2208
rect -5073 1432 -5039 2208
rect -4915 1432 -4881 2208
rect -4757 1432 -4723 2208
rect -4599 1432 -4565 2208
rect -4441 1432 -4407 2208
rect -4283 1432 -4249 2208
rect -4125 1432 -4091 2208
rect -3967 1432 -3933 2208
rect -3809 1432 -3775 2208
rect -3651 1432 -3617 2208
rect -3493 1432 -3459 2208
rect -3335 1432 -3301 2208
rect -3177 1432 -3143 2208
rect -3019 1432 -2985 2208
rect -2861 1432 -2827 2208
rect -2703 1432 -2669 2208
rect -2545 1432 -2511 2208
rect -2387 1432 -2353 2208
rect -2229 1432 -2195 2208
rect -2071 1432 -2037 2208
rect -1913 1432 -1879 2208
rect -1755 1432 -1721 2208
rect -1597 1432 -1563 2208
rect -1439 1432 -1405 2208
rect -1281 1432 -1247 2208
rect -1123 1432 -1089 2208
rect -965 1432 -931 2208
rect -807 1432 -773 2208
rect -649 1432 -615 2208
rect -491 1432 -457 2208
rect -333 1432 -299 2208
rect -175 1432 -141 2208
rect -17 1432 17 2208
rect 141 1432 175 2208
rect 299 1432 333 2208
rect 457 1432 491 2208
rect 615 1432 649 2208
rect 773 1432 807 2208
rect 931 1432 965 2208
rect 1089 1432 1123 2208
rect 1247 1432 1281 2208
rect 1405 1432 1439 2208
rect 1563 1432 1597 2208
rect 1721 1432 1755 2208
rect 1879 1432 1913 2208
rect 2037 1432 2071 2208
rect 2195 1432 2229 2208
rect 2353 1432 2387 2208
rect 2511 1432 2545 2208
rect 2669 1432 2703 2208
rect 2827 1432 2861 2208
rect 2985 1432 3019 2208
rect 3143 1432 3177 2208
rect 3301 1432 3335 2208
rect 3459 1432 3493 2208
rect 3617 1432 3651 2208
rect 3775 1432 3809 2208
rect 3933 1432 3967 2208
rect 4091 1432 4125 2208
rect 4249 1432 4283 2208
rect 4407 1432 4441 2208
rect 4565 1432 4599 2208
rect 4723 1432 4757 2208
rect 4881 1432 4915 2208
rect 5039 1432 5073 2208
rect 5197 1432 5231 2208
rect 5355 1432 5389 2208
rect 5513 1432 5547 2208
rect 5671 1432 5705 2208
rect 5829 1432 5863 2208
rect 5987 1432 6021 2208
rect 6145 1432 6179 2208
rect 6303 1432 6337 2208
rect -6337 522 -6303 1298
rect -6179 522 -6145 1298
rect -6021 522 -5987 1298
rect -5863 522 -5829 1298
rect -5705 522 -5671 1298
rect -5547 522 -5513 1298
rect -5389 522 -5355 1298
rect -5231 522 -5197 1298
rect -5073 522 -5039 1298
rect -4915 522 -4881 1298
rect -4757 522 -4723 1298
rect -4599 522 -4565 1298
rect -4441 522 -4407 1298
rect -4283 522 -4249 1298
rect -4125 522 -4091 1298
rect -3967 522 -3933 1298
rect -3809 522 -3775 1298
rect -3651 522 -3617 1298
rect -3493 522 -3459 1298
rect -3335 522 -3301 1298
rect -3177 522 -3143 1298
rect -3019 522 -2985 1298
rect -2861 522 -2827 1298
rect -2703 522 -2669 1298
rect -2545 522 -2511 1298
rect -2387 522 -2353 1298
rect -2229 522 -2195 1298
rect -2071 522 -2037 1298
rect -1913 522 -1879 1298
rect -1755 522 -1721 1298
rect -1597 522 -1563 1298
rect -1439 522 -1405 1298
rect -1281 522 -1247 1298
rect -1123 522 -1089 1298
rect -965 522 -931 1298
rect -807 522 -773 1298
rect -649 522 -615 1298
rect -491 522 -457 1298
rect -333 522 -299 1298
rect -175 522 -141 1298
rect -17 522 17 1298
rect 141 522 175 1298
rect 299 522 333 1298
rect 457 522 491 1298
rect 615 522 649 1298
rect 773 522 807 1298
rect 931 522 965 1298
rect 1089 522 1123 1298
rect 1247 522 1281 1298
rect 1405 522 1439 1298
rect 1563 522 1597 1298
rect 1721 522 1755 1298
rect 1879 522 1913 1298
rect 2037 522 2071 1298
rect 2195 522 2229 1298
rect 2353 522 2387 1298
rect 2511 522 2545 1298
rect 2669 522 2703 1298
rect 2827 522 2861 1298
rect 2985 522 3019 1298
rect 3143 522 3177 1298
rect 3301 522 3335 1298
rect 3459 522 3493 1298
rect 3617 522 3651 1298
rect 3775 522 3809 1298
rect 3933 522 3967 1298
rect 4091 522 4125 1298
rect 4249 522 4283 1298
rect 4407 522 4441 1298
rect 4565 522 4599 1298
rect 4723 522 4757 1298
rect 4881 522 4915 1298
rect 5039 522 5073 1298
rect 5197 522 5231 1298
rect 5355 522 5389 1298
rect 5513 522 5547 1298
rect 5671 522 5705 1298
rect 5829 522 5863 1298
rect 5987 522 6021 1298
rect 6145 522 6179 1298
rect 6303 522 6337 1298
rect -6337 -388 -6303 388
rect -6179 -388 -6145 388
rect -6021 -388 -5987 388
rect -5863 -388 -5829 388
rect -5705 -388 -5671 388
rect -5547 -388 -5513 388
rect -5389 -388 -5355 388
rect -5231 -388 -5197 388
rect -5073 -388 -5039 388
rect -4915 -388 -4881 388
rect -4757 -388 -4723 388
rect -4599 -388 -4565 388
rect -4441 -388 -4407 388
rect -4283 -388 -4249 388
rect -4125 -388 -4091 388
rect -3967 -388 -3933 388
rect -3809 -388 -3775 388
rect -3651 -388 -3617 388
rect -3493 -388 -3459 388
rect -3335 -388 -3301 388
rect -3177 -388 -3143 388
rect -3019 -388 -2985 388
rect -2861 -388 -2827 388
rect -2703 -388 -2669 388
rect -2545 -388 -2511 388
rect -2387 -388 -2353 388
rect -2229 -388 -2195 388
rect -2071 -388 -2037 388
rect -1913 -388 -1879 388
rect -1755 -388 -1721 388
rect -1597 -388 -1563 388
rect -1439 -388 -1405 388
rect -1281 -388 -1247 388
rect -1123 -388 -1089 388
rect -965 -388 -931 388
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
rect 931 -388 965 388
rect 1089 -388 1123 388
rect 1247 -388 1281 388
rect 1405 -388 1439 388
rect 1563 -388 1597 388
rect 1721 -388 1755 388
rect 1879 -388 1913 388
rect 2037 -388 2071 388
rect 2195 -388 2229 388
rect 2353 -388 2387 388
rect 2511 -388 2545 388
rect 2669 -388 2703 388
rect 2827 -388 2861 388
rect 2985 -388 3019 388
rect 3143 -388 3177 388
rect 3301 -388 3335 388
rect 3459 -388 3493 388
rect 3617 -388 3651 388
rect 3775 -388 3809 388
rect 3933 -388 3967 388
rect 4091 -388 4125 388
rect 4249 -388 4283 388
rect 4407 -388 4441 388
rect 4565 -388 4599 388
rect 4723 -388 4757 388
rect 4881 -388 4915 388
rect 5039 -388 5073 388
rect 5197 -388 5231 388
rect 5355 -388 5389 388
rect 5513 -388 5547 388
rect 5671 -388 5705 388
rect 5829 -388 5863 388
rect 5987 -388 6021 388
rect 6145 -388 6179 388
rect 6303 -388 6337 388
rect -6337 -1298 -6303 -522
rect -6179 -1298 -6145 -522
rect -6021 -1298 -5987 -522
rect -5863 -1298 -5829 -522
rect -5705 -1298 -5671 -522
rect -5547 -1298 -5513 -522
rect -5389 -1298 -5355 -522
rect -5231 -1298 -5197 -522
rect -5073 -1298 -5039 -522
rect -4915 -1298 -4881 -522
rect -4757 -1298 -4723 -522
rect -4599 -1298 -4565 -522
rect -4441 -1298 -4407 -522
rect -4283 -1298 -4249 -522
rect -4125 -1298 -4091 -522
rect -3967 -1298 -3933 -522
rect -3809 -1298 -3775 -522
rect -3651 -1298 -3617 -522
rect -3493 -1298 -3459 -522
rect -3335 -1298 -3301 -522
rect -3177 -1298 -3143 -522
rect -3019 -1298 -2985 -522
rect -2861 -1298 -2827 -522
rect -2703 -1298 -2669 -522
rect -2545 -1298 -2511 -522
rect -2387 -1298 -2353 -522
rect -2229 -1298 -2195 -522
rect -2071 -1298 -2037 -522
rect -1913 -1298 -1879 -522
rect -1755 -1298 -1721 -522
rect -1597 -1298 -1563 -522
rect -1439 -1298 -1405 -522
rect -1281 -1298 -1247 -522
rect -1123 -1298 -1089 -522
rect -965 -1298 -931 -522
rect -807 -1298 -773 -522
rect -649 -1298 -615 -522
rect -491 -1298 -457 -522
rect -333 -1298 -299 -522
rect -175 -1298 -141 -522
rect -17 -1298 17 -522
rect 141 -1298 175 -522
rect 299 -1298 333 -522
rect 457 -1298 491 -522
rect 615 -1298 649 -522
rect 773 -1298 807 -522
rect 931 -1298 965 -522
rect 1089 -1298 1123 -522
rect 1247 -1298 1281 -522
rect 1405 -1298 1439 -522
rect 1563 -1298 1597 -522
rect 1721 -1298 1755 -522
rect 1879 -1298 1913 -522
rect 2037 -1298 2071 -522
rect 2195 -1298 2229 -522
rect 2353 -1298 2387 -522
rect 2511 -1298 2545 -522
rect 2669 -1298 2703 -522
rect 2827 -1298 2861 -522
rect 2985 -1298 3019 -522
rect 3143 -1298 3177 -522
rect 3301 -1298 3335 -522
rect 3459 -1298 3493 -522
rect 3617 -1298 3651 -522
rect 3775 -1298 3809 -522
rect 3933 -1298 3967 -522
rect 4091 -1298 4125 -522
rect 4249 -1298 4283 -522
rect 4407 -1298 4441 -522
rect 4565 -1298 4599 -522
rect 4723 -1298 4757 -522
rect 4881 -1298 4915 -522
rect 5039 -1298 5073 -522
rect 5197 -1298 5231 -522
rect 5355 -1298 5389 -522
rect 5513 -1298 5547 -522
rect 5671 -1298 5705 -522
rect 5829 -1298 5863 -522
rect 5987 -1298 6021 -522
rect 6145 -1298 6179 -522
rect 6303 -1298 6337 -522
rect -6337 -2208 -6303 -1432
rect -6179 -2208 -6145 -1432
rect -6021 -2208 -5987 -1432
rect -5863 -2208 -5829 -1432
rect -5705 -2208 -5671 -1432
rect -5547 -2208 -5513 -1432
rect -5389 -2208 -5355 -1432
rect -5231 -2208 -5197 -1432
rect -5073 -2208 -5039 -1432
rect -4915 -2208 -4881 -1432
rect -4757 -2208 -4723 -1432
rect -4599 -2208 -4565 -1432
rect -4441 -2208 -4407 -1432
rect -4283 -2208 -4249 -1432
rect -4125 -2208 -4091 -1432
rect -3967 -2208 -3933 -1432
rect -3809 -2208 -3775 -1432
rect -3651 -2208 -3617 -1432
rect -3493 -2208 -3459 -1432
rect -3335 -2208 -3301 -1432
rect -3177 -2208 -3143 -1432
rect -3019 -2208 -2985 -1432
rect -2861 -2208 -2827 -1432
rect -2703 -2208 -2669 -1432
rect -2545 -2208 -2511 -1432
rect -2387 -2208 -2353 -1432
rect -2229 -2208 -2195 -1432
rect -2071 -2208 -2037 -1432
rect -1913 -2208 -1879 -1432
rect -1755 -2208 -1721 -1432
rect -1597 -2208 -1563 -1432
rect -1439 -2208 -1405 -1432
rect -1281 -2208 -1247 -1432
rect -1123 -2208 -1089 -1432
rect -965 -2208 -931 -1432
rect -807 -2208 -773 -1432
rect -649 -2208 -615 -1432
rect -491 -2208 -457 -1432
rect -333 -2208 -299 -1432
rect -175 -2208 -141 -1432
rect -17 -2208 17 -1432
rect 141 -2208 175 -1432
rect 299 -2208 333 -1432
rect 457 -2208 491 -1432
rect 615 -2208 649 -1432
rect 773 -2208 807 -1432
rect 931 -2208 965 -1432
rect 1089 -2208 1123 -1432
rect 1247 -2208 1281 -1432
rect 1405 -2208 1439 -1432
rect 1563 -2208 1597 -1432
rect 1721 -2208 1755 -1432
rect 1879 -2208 1913 -1432
rect 2037 -2208 2071 -1432
rect 2195 -2208 2229 -1432
rect 2353 -2208 2387 -1432
rect 2511 -2208 2545 -1432
rect 2669 -2208 2703 -1432
rect 2827 -2208 2861 -1432
rect 2985 -2208 3019 -1432
rect 3143 -2208 3177 -1432
rect 3301 -2208 3335 -1432
rect 3459 -2208 3493 -1432
rect 3617 -2208 3651 -1432
rect 3775 -2208 3809 -1432
rect 3933 -2208 3967 -1432
rect 4091 -2208 4125 -1432
rect 4249 -2208 4283 -1432
rect 4407 -2208 4441 -1432
rect 4565 -2208 4599 -1432
rect 4723 -2208 4757 -1432
rect 4881 -2208 4915 -1432
rect 5039 -2208 5073 -1432
rect 5197 -2208 5231 -1432
rect 5355 -2208 5389 -1432
rect 5513 -2208 5547 -1432
rect 5671 -2208 5705 -1432
rect 5829 -2208 5863 -1432
rect 5987 -2208 6021 -1432
rect 6145 -2208 6179 -1432
rect 6303 -2208 6337 -1432
<< mvpsubdiff >>
rect -6483 2430 6483 2442
rect -6483 2396 -6375 2430
rect 6375 2396 6483 2430
rect -6483 2384 6483 2396
rect -6483 2334 -6425 2384
rect -6483 -2334 -6471 2334
rect -6437 -2334 -6425 2334
rect 6425 2334 6483 2384
rect -6483 -2384 -6425 -2334
rect 6425 -2334 6437 2334
rect 6471 -2334 6483 2334
rect 6425 -2384 6483 -2334
rect -6483 -2396 6483 -2384
rect -6483 -2430 -6375 -2396
rect 6375 -2430 6483 -2396
rect -6483 -2442 6483 -2430
<< mvpsubdiffcont >>
rect -6375 2396 6375 2430
rect -6471 -2334 -6437 2334
rect 6437 -2334 6471 2334
rect -6375 -2430 6375 -2396
<< poly >>
rect -6291 2292 -6191 2308
rect -6291 2258 -6275 2292
rect -6207 2258 -6191 2292
rect -6291 2220 -6191 2258
rect -6133 2292 -6033 2308
rect -6133 2258 -6117 2292
rect -6049 2258 -6033 2292
rect -6133 2220 -6033 2258
rect -5975 2292 -5875 2308
rect -5975 2258 -5959 2292
rect -5891 2258 -5875 2292
rect -5975 2220 -5875 2258
rect -5817 2292 -5717 2308
rect -5817 2258 -5801 2292
rect -5733 2258 -5717 2292
rect -5817 2220 -5717 2258
rect -5659 2292 -5559 2308
rect -5659 2258 -5643 2292
rect -5575 2258 -5559 2292
rect -5659 2220 -5559 2258
rect -5501 2292 -5401 2308
rect -5501 2258 -5485 2292
rect -5417 2258 -5401 2292
rect -5501 2220 -5401 2258
rect -5343 2292 -5243 2308
rect -5343 2258 -5327 2292
rect -5259 2258 -5243 2292
rect -5343 2220 -5243 2258
rect -5185 2292 -5085 2308
rect -5185 2258 -5169 2292
rect -5101 2258 -5085 2292
rect -5185 2220 -5085 2258
rect -5027 2292 -4927 2308
rect -5027 2258 -5011 2292
rect -4943 2258 -4927 2292
rect -5027 2220 -4927 2258
rect -4869 2292 -4769 2308
rect -4869 2258 -4853 2292
rect -4785 2258 -4769 2292
rect -4869 2220 -4769 2258
rect -4711 2292 -4611 2308
rect -4711 2258 -4695 2292
rect -4627 2258 -4611 2292
rect -4711 2220 -4611 2258
rect -4553 2292 -4453 2308
rect -4553 2258 -4537 2292
rect -4469 2258 -4453 2292
rect -4553 2220 -4453 2258
rect -4395 2292 -4295 2308
rect -4395 2258 -4379 2292
rect -4311 2258 -4295 2292
rect -4395 2220 -4295 2258
rect -4237 2292 -4137 2308
rect -4237 2258 -4221 2292
rect -4153 2258 -4137 2292
rect -4237 2220 -4137 2258
rect -4079 2292 -3979 2308
rect -4079 2258 -4063 2292
rect -3995 2258 -3979 2292
rect -4079 2220 -3979 2258
rect -3921 2292 -3821 2308
rect -3921 2258 -3905 2292
rect -3837 2258 -3821 2292
rect -3921 2220 -3821 2258
rect -3763 2292 -3663 2308
rect -3763 2258 -3747 2292
rect -3679 2258 -3663 2292
rect -3763 2220 -3663 2258
rect -3605 2292 -3505 2308
rect -3605 2258 -3589 2292
rect -3521 2258 -3505 2292
rect -3605 2220 -3505 2258
rect -3447 2292 -3347 2308
rect -3447 2258 -3431 2292
rect -3363 2258 -3347 2292
rect -3447 2220 -3347 2258
rect -3289 2292 -3189 2308
rect -3289 2258 -3273 2292
rect -3205 2258 -3189 2292
rect -3289 2220 -3189 2258
rect -3131 2292 -3031 2308
rect -3131 2258 -3115 2292
rect -3047 2258 -3031 2292
rect -3131 2220 -3031 2258
rect -2973 2292 -2873 2308
rect -2973 2258 -2957 2292
rect -2889 2258 -2873 2292
rect -2973 2220 -2873 2258
rect -2815 2292 -2715 2308
rect -2815 2258 -2799 2292
rect -2731 2258 -2715 2292
rect -2815 2220 -2715 2258
rect -2657 2292 -2557 2308
rect -2657 2258 -2641 2292
rect -2573 2258 -2557 2292
rect -2657 2220 -2557 2258
rect -2499 2292 -2399 2308
rect -2499 2258 -2483 2292
rect -2415 2258 -2399 2292
rect -2499 2220 -2399 2258
rect -2341 2292 -2241 2308
rect -2341 2258 -2325 2292
rect -2257 2258 -2241 2292
rect -2341 2220 -2241 2258
rect -2183 2292 -2083 2308
rect -2183 2258 -2167 2292
rect -2099 2258 -2083 2292
rect -2183 2220 -2083 2258
rect -2025 2292 -1925 2308
rect -2025 2258 -2009 2292
rect -1941 2258 -1925 2292
rect -2025 2220 -1925 2258
rect -1867 2292 -1767 2308
rect -1867 2258 -1851 2292
rect -1783 2258 -1767 2292
rect -1867 2220 -1767 2258
rect -1709 2292 -1609 2308
rect -1709 2258 -1693 2292
rect -1625 2258 -1609 2292
rect -1709 2220 -1609 2258
rect -1551 2292 -1451 2308
rect -1551 2258 -1535 2292
rect -1467 2258 -1451 2292
rect -1551 2220 -1451 2258
rect -1393 2292 -1293 2308
rect -1393 2258 -1377 2292
rect -1309 2258 -1293 2292
rect -1393 2220 -1293 2258
rect -1235 2292 -1135 2308
rect -1235 2258 -1219 2292
rect -1151 2258 -1135 2292
rect -1235 2220 -1135 2258
rect -1077 2292 -977 2308
rect -1077 2258 -1061 2292
rect -993 2258 -977 2292
rect -1077 2220 -977 2258
rect -919 2292 -819 2308
rect -919 2258 -903 2292
rect -835 2258 -819 2292
rect -919 2220 -819 2258
rect -761 2292 -661 2308
rect -761 2258 -745 2292
rect -677 2258 -661 2292
rect -761 2220 -661 2258
rect -603 2292 -503 2308
rect -603 2258 -587 2292
rect -519 2258 -503 2292
rect -603 2220 -503 2258
rect -445 2292 -345 2308
rect -445 2258 -429 2292
rect -361 2258 -345 2292
rect -445 2220 -345 2258
rect -287 2292 -187 2308
rect -287 2258 -271 2292
rect -203 2258 -187 2292
rect -287 2220 -187 2258
rect -129 2292 -29 2308
rect -129 2258 -113 2292
rect -45 2258 -29 2292
rect -129 2220 -29 2258
rect 29 2292 129 2308
rect 29 2258 45 2292
rect 113 2258 129 2292
rect 29 2220 129 2258
rect 187 2292 287 2308
rect 187 2258 203 2292
rect 271 2258 287 2292
rect 187 2220 287 2258
rect 345 2292 445 2308
rect 345 2258 361 2292
rect 429 2258 445 2292
rect 345 2220 445 2258
rect 503 2292 603 2308
rect 503 2258 519 2292
rect 587 2258 603 2292
rect 503 2220 603 2258
rect 661 2292 761 2308
rect 661 2258 677 2292
rect 745 2258 761 2292
rect 661 2220 761 2258
rect 819 2292 919 2308
rect 819 2258 835 2292
rect 903 2258 919 2292
rect 819 2220 919 2258
rect 977 2292 1077 2308
rect 977 2258 993 2292
rect 1061 2258 1077 2292
rect 977 2220 1077 2258
rect 1135 2292 1235 2308
rect 1135 2258 1151 2292
rect 1219 2258 1235 2292
rect 1135 2220 1235 2258
rect 1293 2292 1393 2308
rect 1293 2258 1309 2292
rect 1377 2258 1393 2292
rect 1293 2220 1393 2258
rect 1451 2292 1551 2308
rect 1451 2258 1467 2292
rect 1535 2258 1551 2292
rect 1451 2220 1551 2258
rect 1609 2292 1709 2308
rect 1609 2258 1625 2292
rect 1693 2258 1709 2292
rect 1609 2220 1709 2258
rect 1767 2292 1867 2308
rect 1767 2258 1783 2292
rect 1851 2258 1867 2292
rect 1767 2220 1867 2258
rect 1925 2292 2025 2308
rect 1925 2258 1941 2292
rect 2009 2258 2025 2292
rect 1925 2220 2025 2258
rect 2083 2292 2183 2308
rect 2083 2258 2099 2292
rect 2167 2258 2183 2292
rect 2083 2220 2183 2258
rect 2241 2292 2341 2308
rect 2241 2258 2257 2292
rect 2325 2258 2341 2292
rect 2241 2220 2341 2258
rect 2399 2292 2499 2308
rect 2399 2258 2415 2292
rect 2483 2258 2499 2292
rect 2399 2220 2499 2258
rect 2557 2292 2657 2308
rect 2557 2258 2573 2292
rect 2641 2258 2657 2292
rect 2557 2220 2657 2258
rect 2715 2292 2815 2308
rect 2715 2258 2731 2292
rect 2799 2258 2815 2292
rect 2715 2220 2815 2258
rect 2873 2292 2973 2308
rect 2873 2258 2889 2292
rect 2957 2258 2973 2292
rect 2873 2220 2973 2258
rect 3031 2292 3131 2308
rect 3031 2258 3047 2292
rect 3115 2258 3131 2292
rect 3031 2220 3131 2258
rect 3189 2292 3289 2308
rect 3189 2258 3205 2292
rect 3273 2258 3289 2292
rect 3189 2220 3289 2258
rect 3347 2292 3447 2308
rect 3347 2258 3363 2292
rect 3431 2258 3447 2292
rect 3347 2220 3447 2258
rect 3505 2292 3605 2308
rect 3505 2258 3521 2292
rect 3589 2258 3605 2292
rect 3505 2220 3605 2258
rect 3663 2292 3763 2308
rect 3663 2258 3679 2292
rect 3747 2258 3763 2292
rect 3663 2220 3763 2258
rect 3821 2292 3921 2308
rect 3821 2258 3837 2292
rect 3905 2258 3921 2292
rect 3821 2220 3921 2258
rect 3979 2292 4079 2308
rect 3979 2258 3995 2292
rect 4063 2258 4079 2292
rect 3979 2220 4079 2258
rect 4137 2292 4237 2308
rect 4137 2258 4153 2292
rect 4221 2258 4237 2292
rect 4137 2220 4237 2258
rect 4295 2292 4395 2308
rect 4295 2258 4311 2292
rect 4379 2258 4395 2292
rect 4295 2220 4395 2258
rect 4453 2292 4553 2308
rect 4453 2258 4469 2292
rect 4537 2258 4553 2292
rect 4453 2220 4553 2258
rect 4611 2292 4711 2308
rect 4611 2258 4627 2292
rect 4695 2258 4711 2292
rect 4611 2220 4711 2258
rect 4769 2292 4869 2308
rect 4769 2258 4785 2292
rect 4853 2258 4869 2292
rect 4769 2220 4869 2258
rect 4927 2292 5027 2308
rect 4927 2258 4943 2292
rect 5011 2258 5027 2292
rect 4927 2220 5027 2258
rect 5085 2292 5185 2308
rect 5085 2258 5101 2292
rect 5169 2258 5185 2292
rect 5085 2220 5185 2258
rect 5243 2292 5343 2308
rect 5243 2258 5259 2292
rect 5327 2258 5343 2292
rect 5243 2220 5343 2258
rect 5401 2292 5501 2308
rect 5401 2258 5417 2292
rect 5485 2258 5501 2292
rect 5401 2220 5501 2258
rect 5559 2292 5659 2308
rect 5559 2258 5575 2292
rect 5643 2258 5659 2292
rect 5559 2220 5659 2258
rect 5717 2292 5817 2308
rect 5717 2258 5733 2292
rect 5801 2258 5817 2292
rect 5717 2220 5817 2258
rect 5875 2292 5975 2308
rect 5875 2258 5891 2292
rect 5959 2258 5975 2292
rect 5875 2220 5975 2258
rect 6033 2292 6133 2308
rect 6033 2258 6049 2292
rect 6117 2258 6133 2292
rect 6033 2220 6133 2258
rect 6191 2292 6291 2308
rect 6191 2258 6207 2292
rect 6275 2258 6291 2292
rect 6191 2220 6291 2258
rect -6291 1382 -6191 1420
rect -6291 1348 -6275 1382
rect -6207 1348 -6191 1382
rect -6291 1310 -6191 1348
rect -6133 1382 -6033 1420
rect -6133 1348 -6117 1382
rect -6049 1348 -6033 1382
rect -6133 1310 -6033 1348
rect -5975 1382 -5875 1420
rect -5975 1348 -5959 1382
rect -5891 1348 -5875 1382
rect -5975 1310 -5875 1348
rect -5817 1382 -5717 1420
rect -5817 1348 -5801 1382
rect -5733 1348 -5717 1382
rect -5817 1310 -5717 1348
rect -5659 1382 -5559 1420
rect -5659 1348 -5643 1382
rect -5575 1348 -5559 1382
rect -5659 1310 -5559 1348
rect -5501 1382 -5401 1420
rect -5501 1348 -5485 1382
rect -5417 1348 -5401 1382
rect -5501 1310 -5401 1348
rect -5343 1382 -5243 1420
rect -5343 1348 -5327 1382
rect -5259 1348 -5243 1382
rect -5343 1310 -5243 1348
rect -5185 1382 -5085 1420
rect -5185 1348 -5169 1382
rect -5101 1348 -5085 1382
rect -5185 1310 -5085 1348
rect -5027 1382 -4927 1420
rect -5027 1348 -5011 1382
rect -4943 1348 -4927 1382
rect -5027 1310 -4927 1348
rect -4869 1382 -4769 1420
rect -4869 1348 -4853 1382
rect -4785 1348 -4769 1382
rect -4869 1310 -4769 1348
rect -4711 1382 -4611 1420
rect -4711 1348 -4695 1382
rect -4627 1348 -4611 1382
rect -4711 1310 -4611 1348
rect -4553 1382 -4453 1420
rect -4553 1348 -4537 1382
rect -4469 1348 -4453 1382
rect -4553 1310 -4453 1348
rect -4395 1382 -4295 1420
rect -4395 1348 -4379 1382
rect -4311 1348 -4295 1382
rect -4395 1310 -4295 1348
rect -4237 1382 -4137 1420
rect -4237 1348 -4221 1382
rect -4153 1348 -4137 1382
rect -4237 1310 -4137 1348
rect -4079 1382 -3979 1420
rect -4079 1348 -4063 1382
rect -3995 1348 -3979 1382
rect -4079 1310 -3979 1348
rect -3921 1382 -3821 1420
rect -3921 1348 -3905 1382
rect -3837 1348 -3821 1382
rect -3921 1310 -3821 1348
rect -3763 1382 -3663 1420
rect -3763 1348 -3747 1382
rect -3679 1348 -3663 1382
rect -3763 1310 -3663 1348
rect -3605 1382 -3505 1420
rect -3605 1348 -3589 1382
rect -3521 1348 -3505 1382
rect -3605 1310 -3505 1348
rect -3447 1382 -3347 1420
rect -3447 1348 -3431 1382
rect -3363 1348 -3347 1382
rect -3447 1310 -3347 1348
rect -3289 1382 -3189 1420
rect -3289 1348 -3273 1382
rect -3205 1348 -3189 1382
rect -3289 1310 -3189 1348
rect -3131 1382 -3031 1420
rect -3131 1348 -3115 1382
rect -3047 1348 -3031 1382
rect -3131 1310 -3031 1348
rect -2973 1382 -2873 1420
rect -2973 1348 -2957 1382
rect -2889 1348 -2873 1382
rect -2973 1310 -2873 1348
rect -2815 1382 -2715 1420
rect -2815 1348 -2799 1382
rect -2731 1348 -2715 1382
rect -2815 1310 -2715 1348
rect -2657 1382 -2557 1420
rect -2657 1348 -2641 1382
rect -2573 1348 -2557 1382
rect -2657 1310 -2557 1348
rect -2499 1382 -2399 1420
rect -2499 1348 -2483 1382
rect -2415 1348 -2399 1382
rect -2499 1310 -2399 1348
rect -2341 1382 -2241 1420
rect -2341 1348 -2325 1382
rect -2257 1348 -2241 1382
rect -2341 1310 -2241 1348
rect -2183 1382 -2083 1420
rect -2183 1348 -2167 1382
rect -2099 1348 -2083 1382
rect -2183 1310 -2083 1348
rect -2025 1382 -1925 1420
rect -2025 1348 -2009 1382
rect -1941 1348 -1925 1382
rect -2025 1310 -1925 1348
rect -1867 1382 -1767 1420
rect -1867 1348 -1851 1382
rect -1783 1348 -1767 1382
rect -1867 1310 -1767 1348
rect -1709 1382 -1609 1420
rect -1709 1348 -1693 1382
rect -1625 1348 -1609 1382
rect -1709 1310 -1609 1348
rect -1551 1382 -1451 1420
rect -1551 1348 -1535 1382
rect -1467 1348 -1451 1382
rect -1551 1310 -1451 1348
rect -1393 1382 -1293 1420
rect -1393 1348 -1377 1382
rect -1309 1348 -1293 1382
rect -1393 1310 -1293 1348
rect -1235 1382 -1135 1420
rect -1235 1348 -1219 1382
rect -1151 1348 -1135 1382
rect -1235 1310 -1135 1348
rect -1077 1382 -977 1420
rect -1077 1348 -1061 1382
rect -993 1348 -977 1382
rect -1077 1310 -977 1348
rect -919 1382 -819 1420
rect -919 1348 -903 1382
rect -835 1348 -819 1382
rect -919 1310 -819 1348
rect -761 1382 -661 1420
rect -761 1348 -745 1382
rect -677 1348 -661 1382
rect -761 1310 -661 1348
rect -603 1382 -503 1420
rect -603 1348 -587 1382
rect -519 1348 -503 1382
rect -603 1310 -503 1348
rect -445 1382 -345 1420
rect -445 1348 -429 1382
rect -361 1348 -345 1382
rect -445 1310 -345 1348
rect -287 1382 -187 1420
rect -287 1348 -271 1382
rect -203 1348 -187 1382
rect -287 1310 -187 1348
rect -129 1382 -29 1420
rect -129 1348 -113 1382
rect -45 1348 -29 1382
rect -129 1310 -29 1348
rect 29 1382 129 1420
rect 29 1348 45 1382
rect 113 1348 129 1382
rect 29 1310 129 1348
rect 187 1382 287 1420
rect 187 1348 203 1382
rect 271 1348 287 1382
rect 187 1310 287 1348
rect 345 1382 445 1420
rect 345 1348 361 1382
rect 429 1348 445 1382
rect 345 1310 445 1348
rect 503 1382 603 1420
rect 503 1348 519 1382
rect 587 1348 603 1382
rect 503 1310 603 1348
rect 661 1382 761 1420
rect 661 1348 677 1382
rect 745 1348 761 1382
rect 661 1310 761 1348
rect 819 1382 919 1420
rect 819 1348 835 1382
rect 903 1348 919 1382
rect 819 1310 919 1348
rect 977 1382 1077 1420
rect 977 1348 993 1382
rect 1061 1348 1077 1382
rect 977 1310 1077 1348
rect 1135 1382 1235 1420
rect 1135 1348 1151 1382
rect 1219 1348 1235 1382
rect 1135 1310 1235 1348
rect 1293 1382 1393 1420
rect 1293 1348 1309 1382
rect 1377 1348 1393 1382
rect 1293 1310 1393 1348
rect 1451 1382 1551 1420
rect 1451 1348 1467 1382
rect 1535 1348 1551 1382
rect 1451 1310 1551 1348
rect 1609 1382 1709 1420
rect 1609 1348 1625 1382
rect 1693 1348 1709 1382
rect 1609 1310 1709 1348
rect 1767 1382 1867 1420
rect 1767 1348 1783 1382
rect 1851 1348 1867 1382
rect 1767 1310 1867 1348
rect 1925 1382 2025 1420
rect 1925 1348 1941 1382
rect 2009 1348 2025 1382
rect 1925 1310 2025 1348
rect 2083 1382 2183 1420
rect 2083 1348 2099 1382
rect 2167 1348 2183 1382
rect 2083 1310 2183 1348
rect 2241 1382 2341 1420
rect 2241 1348 2257 1382
rect 2325 1348 2341 1382
rect 2241 1310 2341 1348
rect 2399 1382 2499 1420
rect 2399 1348 2415 1382
rect 2483 1348 2499 1382
rect 2399 1310 2499 1348
rect 2557 1382 2657 1420
rect 2557 1348 2573 1382
rect 2641 1348 2657 1382
rect 2557 1310 2657 1348
rect 2715 1382 2815 1420
rect 2715 1348 2731 1382
rect 2799 1348 2815 1382
rect 2715 1310 2815 1348
rect 2873 1382 2973 1420
rect 2873 1348 2889 1382
rect 2957 1348 2973 1382
rect 2873 1310 2973 1348
rect 3031 1382 3131 1420
rect 3031 1348 3047 1382
rect 3115 1348 3131 1382
rect 3031 1310 3131 1348
rect 3189 1382 3289 1420
rect 3189 1348 3205 1382
rect 3273 1348 3289 1382
rect 3189 1310 3289 1348
rect 3347 1382 3447 1420
rect 3347 1348 3363 1382
rect 3431 1348 3447 1382
rect 3347 1310 3447 1348
rect 3505 1382 3605 1420
rect 3505 1348 3521 1382
rect 3589 1348 3605 1382
rect 3505 1310 3605 1348
rect 3663 1382 3763 1420
rect 3663 1348 3679 1382
rect 3747 1348 3763 1382
rect 3663 1310 3763 1348
rect 3821 1382 3921 1420
rect 3821 1348 3837 1382
rect 3905 1348 3921 1382
rect 3821 1310 3921 1348
rect 3979 1382 4079 1420
rect 3979 1348 3995 1382
rect 4063 1348 4079 1382
rect 3979 1310 4079 1348
rect 4137 1382 4237 1420
rect 4137 1348 4153 1382
rect 4221 1348 4237 1382
rect 4137 1310 4237 1348
rect 4295 1382 4395 1420
rect 4295 1348 4311 1382
rect 4379 1348 4395 1382
rect 4295 1310 4395 1348
rect 4453 1382 4553 1420
rect 4453 1348 4469 1382
rect 4537 1348 4553 1382
rect 4453 1310 4553 1348
rect 4611 1382 4711 1420
rect 4611 1348 4627 1382
rect 4695 1348 4711 1382
rect 4611 1310 4711 1348
rect 4769 1382 4869 1420
rect 4769 1348 4785 1382
rect 4853 1348 4869 1382
rect 4769 1310 4869 1348
rect 4927 1382 5027 1420
rect 4927 1348 4943 1382
rect 5011 1348 5027 1382
rect 4927 1310 5027 1348
rect 5085 1382 5185 1420
rect 5085 1348 5101 1382
rect 5169 1348 5185 1382
rect 5085 1310 5185 1348
rect 5243 1382 5343 1420
rect 5243 1348 5259 1382
rect 5327 1348 5343 1382
rect 5243 1310 5343 1348
rect 5401 1382 5501 1420
rect 5401 1348 5417 1382
rect 5485 1348 5501 1382
rect 5401 1310 5501 1348
rect 5559 1382 5659 1420
rect 5559 1348 5575 1382
rect 5643 1348 5659 1382
rect 5559 1310 5659 1348
rect 5717 1382 5817 1420
rect 5717 1348 5733 1382
rect 5801 1348 5817 1382
rect 5717 1310 5817 1348
rect 5875 1382 5975 1420
rect 5875 1348 5891 1382
rect 5959 1348 5975 1382
rect 5875 1310 5975 1348
rect 6033 1382 6133 1420
rect 6033 1348 6049 1382
rect 6117 1348 6133 1382
rect 6033 1310 6133 1348
rect 6191 1382 6291 1420
rect 6191 1348 6207 1382
rect 6275 1348 6291 1382
rect 6191 1310 6291 1348
rect -6291 472 -6191 510
rect -6291 438 -6275 472
rect -6207 438 -6191 472
rect -6291 400 -6191 438
rect -6133 472 -6033 510
rect -6133 438 -6117 472
rect -6049 438 -6033 472
rect -6133 400 -6033 438
rect -5975 472 -5875 510
rect -5975 438 -5959 472
rect -5891 438 -5875 472
rect -5975 400 -5875 438
rect -5817 472 -5717 510
rect -5817 438 -5801 472
rect -5733 438 -5717 472
rect -5817 400 -5717 438
rect -5659 472 -5559 510
rect -5659 438 -5643 472
rect -5575 438 -5559 472
rect -5659 400 -5559 438
rect -5501 472 -5401 510
rect -5501 438 -5485 472
rect -5417 438 -5401 472
rect -5501 400 -5401 438
rect -5343 472 -5243 510
rect -5343 438 -5327 472
rect -5259 438 -5243 472
rect -5343 400 -5243 438
rect -5185 472 -5085 510
rect -5185 438 -5169 472
rect -5101 438 -5085 472
rect -5185 400 -5085 438
rect -5027 472 -4927 510
rect -5027 438 -5011 472
rect -4943 438 -4927 472
rect -5027 400 -4927 438
rect -4869 472 -4769 510
rect -4869 438 -4853 472
rect -4785 438 -4769 472
rect -4869 400 -4769 438
rect -4711 472 -4611 510
rect -4711 438 -4695 472
rect -4627 438 -4611 472
rect -4711 400 -4611 438
rect -4553 472 -4453 510
rect -4553 438 -4537 472
rect -4469 438 -4453 472
rect -4553 400 -4453 438
rect -4395 472 -4295 510
rect -4395 438 -4379 472
rect -4311 438 -4295 472
rect -4395 400 -4295 438
rect -4237 472 -4137 510
rect -4237 438 -4221 472
rect -4153 438 -4137 472
rect -4237 400 -4137 438
rect -4079 472 -3979 510
rect -4079 438 -4063 472
rect -3995 438 -3979 472
rect -4079 400 -3979 438
rect -3921 472 -3821 510
rect -3921 438 -3905 472
rect -3837 438 -3821 472
rect -3921 400 -3821 438
rect -3763 472 -3663 510
rect -3763 438 -3747 472
rect -3679 438 -3663 472
rect -3763 400 -3663 438
rect -3605 472 -3505 510
rect -3605 438 -3589 472
rect -3521 438 -3505 472
rect -3605 400 -3505 438
rect -3447 472 -3347 510
rect -3447 438 -3431 472
rect -3363 438 -3347 472
rect -3447 400 -3347 438
rect -3289 472 -3189 510
rect -3289 438 -3273 472
rect -3205 438 -3189 472
rect -3289 400 -3189 438
rect -3131 472 -3031 510
rect -3131 438 -3115 472
rect -3047 438 -3031 472
rect -3131 400 -3031 438
rect -2973 472 -2873 510
rect -2973 438 -2957 472
rect -2889 438 -2873 472
rect -2973 400 -2873 438
rect -2815 472 -2715 510
rect -2815 438 -2799 472
rect -2731 438 -2715 472
rect -2815 400 -2715 438
rect -2657 472 -2557 510
rect -2657 438 -2641 472
rect -2573 438 -2557 472
rect -2657 400 -2557 438
rect -2499 472 -2399 510
rect -2499 438 -2483 472
rect -2415 438 -2399 472
rect -2499 400 -2399 438
rect -2341 472 -2241 510
rect -2341 438 -2325 472
rect -2257 438 -2241 472
rect -2341 400 -2241 438
rect -2183 472 -2083 510
rect -2183 438 -2167 472
rect -2099 438 -2083 472
rect -2183 400 -2083 438
rect -2025 472 -1925 510
rect -2025 438 -2009 472
rect -1941 438 -1925 472
rect -2025 400 -1925 438
rect -1867 472 -1767 510
rect -1867 438 -1851 472
rect -1783 438 -1767 472
rect -1867 400 -1767 438
rect -1709 472 -1609 510
rect -1709 438 -1693 472
rect -1625 438 -1609 472
rect -1709 400 -1609 438
rect -1551 472 -1451 510
rect -1551 438 -1535 472
rect -1467 438 -1451 472
rect -1551 400 -1451 438
rect -1393 472 -1293 510
rect -1393 438 -1377 472
rect -1309 438 -1293 472
rect -1393 400 -1293 438
rect -1235 472 -1135 510
rect -1235 438 -1219 472
rect -1151 438 -1135 472
rect -1235 400 -1135 438
rect -1077 472 -977 510
rect -1077 438 -1061 472
rect -993 438 -977 472
rect -1077 400 -977 438
rect -919 472 -819 510
rect -919 438 -903 472
rect -835 438 -819 472
rect -919 400 -819 438
rect -761 472 -661 510
rect -761 438 -745 472
rect -677 438 -661 472
rect -761 400 -661 438
rect -603 472 -503 510
rect -603 438 -587 472
rect -519 438 -503 472
rect -603 400 -503 438
rect -445 472 -345 510
rect -445 438 -429 472
rect -361 438 -345 472
rect -445 400 -345 438
rect -287 472 -187 510
rect -287 438 -271 472
rect -203 438 -187 472
rect -287 400 -187 438
rect -129 472 -29 510
rect -129 438 -113 472
rect -45 438 -29 472
rect -129 400 -29 438
rect 29 472 129 510
rect 29 438 45 472
rect 113 438 129 472
rect 29 400 129 438
rect 187 472 287 510
rect 187 438 203 472
rect 271 438 287 472
rect 187 400 287 438
rect 345 472 445 510
rect 345 438 361 472
rect 429 438 445 472
rect 345 400 445 438
rect 503 472 603 510
rect 503 438 519 472
rect 587 438 603 472
rect 503 400 603 438
rect 661 472 761 510
rect 661 438 677 472
rect 745 438 761 472
rect 661 400 761 438
rect 819 472 919 510
rect 819 438 835 472
rect 903 438 919 472
rect 819 400 919 438
rect 977 472 1077 510
rect 977 438 993 472
rect 1061 438 1077 472
rect 977 400 1077 438
rect 1135 472 1235 510
rect 1135 438 1151 472
rect 1219 438 1235 472
rect 1135 400 1235 438
rect 1293 472 1393 510
rect 1293 438 1309 472
rect 1377 438 1393 472
rect 1293 400 1393 438
rect 1451 472 1551 510
rect 1451 438 1467 472
rect 1535 438 1551 472
rect 1451 400 1551 438
rect 1609 472 1709 510
rect 1609 438 1625 472
rect 1693 438 1709 472
rect 1609 400 1709 438
rect 1767 472 1867 510
rect 1767 438 1783 472
rect 1851 438 1867 472
rect 1767 400 1867 438
rect 1925 472 2025 510
rect 1925 438 1941 472
rect 2009 438 2025 472
rect 1925 400 2025 438
rect 2083 472 2183 510
rect 2083 438 2099 472
rect 2167 438 2183 472
rect 2083 400 2183 438
rect 2241 472 2341 510
rect 2241 438 2257 472
rect 2325 438 2341 472
rect 2241 400 2341 438
rect 2399 472 2499 510
rect 2399 438 2415 472
rect 2483 438 2499 472
rect 2399 400 2499 438
rect 2557 472 2657 510
rect 2557 438 2573 472
rect 2641 438 2657 472
rect 2557 400 2657 438
rect 2715 472 2815 510
rect 2715 438 2731 472
rect 2799 438 2815 472
rect 2715 400 2815 438
rect 2873 472 2973 510
rect 2873 438 2889 472
rect 2957 438 2973 472
rect 2873 400 2973 438
rect 3031 472 3131 510
rect 3031 438 3047 472
rect 3115 438 3131 472
rect 3031 400 3131 438
rect 3189 472 3289 510
rect 3189 438 3205 472
rect 3273 438 3289 472
rect 3189 400 3289 438
rect 3347 472 3447 510
rect 3347 438 3363 472
rect 3431 438 3447 472
rect 3347 400 3447 438
rect 3505 472 3605 510
rect 3505 438 3521 472
rect 3589 438 3605 472
rect 3505 400 3605 438
rect 3663 472 3763 510
rect 3663 438 3679 472
rect 3747 438 3763 472
rect 3663 400 3763 438
rect 3821 472 3921 510
rect 3821 438 3837 472
rect 3905 438 3921 472
rect 3821 400 3921 438
rect 3979 472 4079 510
rect 3979 438 3995 472
rect 4063 438 4079 472
rect 3979 400 4079 438
rect 4137 472 4237 510
rect 4137 438 4153 472
rect 4221 438 4237 472
rect 4137 400 4237 438
rect 4295 472 4395 510
rect 4295 438 4311 472
rect 4379 438 4395 472
rect 4295 400 4395 438
rect 4453 472 4553 510
rect 4453 438 4469 472
rect 4537 438 4553 472
rect 4453 400 4553 438
rect 4611 472 4711 510
rect 4611 438 4627 472
rect 4695 438 4711 472
rect 4611 400 4711 438
rect 4769 472 4869 510
rect 4769 438 4785 472
rect 4853 438 4869 472
rect 4769 400 4869 438
rect 4927 472 5027 510
rect 4927 438 4943 472
rect 5011 438 5027 472
rect 4927 400 5027 438
rect 5085 472 5185 510
rect 5085 438 5101 472
rect 5169 438 5185 472
rect 5085 400 5185 438
rect 5243 472 5343 510
rect 5243 438 5259 472
rect 5327 438 5343 472
rect 5243 400 5343 438
rect 5401 472 5501 510
rect 5401 438 5417 472
rect 5485 438 5501 472
rect 5401 400 5501 438
rect 5559 472 5659 510
rect 5559 438 5575 472
rect 5643 438 5659 472
rect 5559 400 5659 438
rect 5717 472 5817 510
rect 5717 438 5733 472
rect 5801 438 5817 472
rect 5717 400 5817 438
rect 5875 472 5975 510
rect 5875 438 5891 472
rect 5959 438 5975 472
rect 5875 400 5975 438
rect 6033 472 6133 510
rect 6033 438 6049 472
rect 6117 438 6133 472
rect 6033 400 6133 438
rect 6191 472 6291 510
rect 6191 438 6207 472
rect 6275 438 6291 472
rect 6191 400 6291 438
rect -6291 -438 -6191 -400
rect -6291 -472 -6275 -438
rect -6207 -472 -6191 -438
rect -6291 -510 -6191 -472
rect -6133 -438 -6033 -400
rect -6133 -472 -6117 -438
rect -6049 -472 -6033 -438
rect -6133 -510 -6033 -472
rect -5975 -438 -5875 -400
rect -5975 -472 -5959 -438
rect -5891 -472 -5875 -438
rect -5975 -510 -5875 -472
rect -5817 -438 -5717 -400
rect -5817 -472 -5801 -438
rect -5733 -472 -5717 -438
rect -5817 -510 -5717 -472
rect -5659 -438 -5559 -400
rect -5659 -472 -5643 -438
rect -5575 -472 -5559 -438
rect -5659 -510 -5559 -472
rect -5501 -438 -5401 -400
rect -5501 -472 -5485 -438
rect -5417 -472 -5401 -438
rect -5501 -510 -5401 -472
rect -5343 -438 -5243 -400
rect -5343 -472 -5327 -438
rect -5259 -472 -5243 -438
rect -5343 -510 -5243 -472
rect -5185 -438 -5085 -400
rect -5185 -472 -5169 -438
rect -5101 -472 -5085 -438
rect -5185 -510 -5085 -472
rect -5027 -438 -4927 -400
rect -5027 -472 -5011 -438
rect -4943 -472 -4927 -438
rect -5027 -510 -4927 -472
rect -4869 -438 -4769 -400
rect -4869 -472 -4853 -438
rect -4785 -472 -4769 -438
rect -4869 -510 -4769 -472
rect -4711 -438 -4611 -400
rect -4711 -472 -4695 -438
rect -4627 -472 -4611 -438
rect -4711 -510 -4611 -472
rect -4553 -438 -4453 -400
rect -4553 -472 -4537 -438
rect -4469 -472 -4453 -438
rect -4553 -510 -4453 -472
rect -4395 -438 -4295 -400
rect -4395 -472 -4379 -438
rect -4311 -472 -4295 -438
rect -4395 -510 -4295 -472
rect -4237 -438 -4137 -400
rect -4237 -472 -4221 -438
rect -4153 -472 -4137 -438
rect -4237 -510 -4137 -472
rect -4079 -438 -3979 -400
rect -4079 -472 -4063 -438
rect -3995 -472 -3979 -438
rect -4079 -510 -3979 -472
rect -3921 -438 -3821 -400
rect -3921 -472 -3905 -438
rect -3837 -472 -3821 -438
rect -3921 -510 -3821 -472
rect -3763 -438 -3663 -400
rect -3763 -472 -3747 -438
rect -3679 -472 -3663 -438
rect -3763 -510 -3663 -472
rect -3605 -438 -3505 -400
rect -3605 -472 -3589 -438
rect -3521 -472 -3505 -438
rect -3605 -510 -3505 -472
rect -3447 -438 -3347 -400
rect -3447 -472 -3431 -438
rect -3363 -472 -3347 -438
rect -3447 -510 -3347 -472
rect -3289 -438 -3189 -400
rect -3289 -472 -3273 -438
rect -3205 -472 -3189 -438
rect -3289 -510 -3189 -472
rect -3131 -438 -3031 -400
rect -3131 -472 -3115 -438
rect -3047 -472 -3031 -438
rect -3131 -510 -3031 -472
rect -2973 -438 -2873 -400
rect -2973 -472 -2957 -438
rect -2889 -472 -2873 -438
rect -2973 -510 -2873 -472
rect -2815 -438 -2715 -400
rect -2815 -472 -2799 -438
rect -2731 -472 -2715 -438
rect -2815 -510 -2715 -472
rect -2657 -438 -2557 -400
rect -2657 -472 -2641 -438
rect -2573 -472 -2557 -438
rect -2657 -510 -2557 -472
rect -2499 -438 -2399 -400
rect -2499 -472 -2483 -438
rect -2415 -472 -2399 -438
rect -2499 -510 -2399 -472
rect -2341 -438 -2241 -400
rect -2341 -472 -2325 -438
rect -2257 -472 -2241 -438
rect -2341 -510 -2241 -472
rect -2183 -438 -2083 -400
rect -2183 -472 -2167 -438
rect -2099 -472 -2083 -438
rect -2183 -510 -2083 -472
rect -2025 -438 -1925 -400
rect -2025 -472 -2009 -438
rect -1941 -472 -1925 -438
rect -2025 -510 -1925 -472
rect -1867 -438 -1767 -400
rect -1867 -472 -1851 -438
rect -1783 -472 -1767 -438
rect -1867 -510 -1767 -472
rect -1709 -438 -1609 -400
rect -1709 -472 -1693 -438
rect -1625 -472 -1609 -438
rect -1709 -510 -1609 -472
rect -1551 -438 -1451 -400
rect -1551 -472 -1535 -438
rect -1467 -472 -1451 -438
rect -1551 -510 -1451 -472
rect -1393 -438 -1293 -400
rect -1393 -472 -1377 -438
rect -1309 -472 -1293 -438
rect -1393 -510 -1293 -472
rect -1235 -438 -1135 -400
rect -1235 -472 -1219 -438
rect -1151 -472 -1135 -438
rect -1235 -510 -1135 -472
rect -1077 -438 -977 -400
rect -1077 -472 -1061 -438
rect -993 -472 -977 -438
rect -1077 -510 -977 -472
rect -919 -438 -819 -400
rect -919 -472 -903 -438
rect -835 -472 -819 -438
rect -919 -510 -819 -472
rect -761 -438 -661 -400
rect -761 -472 -745 -438
rect -677 -472 -661 -438
rect -761 -510 -661 -472
rect -603 -438 -503 -400
rect -603 -472 -587 -438
rect -519 -472 -503 -438
rect -603 -510 -503 -472
rect -445 -438 -345 -400
rect -445 -472 -429 -438
rect -361 -472 -345 -438
rect -445 -510 -345 -472
rect -287 -438 -187 -400
rect -287 -472 -271 -438
rect -203 -472 -187 -438
rect -287 -510 -187 -472
rect -129 -438 -29 -400
rect -129 -472 -113 -438
rect -45 -472 -29 -438
rect -129 -510 -29 -472
rect 29 -438 129 -400
rect 29 -472 45 -438
rect 113 -472 129 -438
rect 29 -510 129 -472
rect 187 -438 287 -400
rect 187 -472 203 -438
rect 271 -472 287 -438
rect 187 -510 287 -472
rect 345 -438 445 -400
rect 345 -472 361 -438
rect 429 -472 445 -438
rect 345 -510 445 -472
rect 503 -438 603 -400
rect 503 -472 519 -438
rect 587 -472 603 -438
rect 503 -510 603 -472
rect 661 -438 761 -400
rect 661 -472 677 -438
rect 745 -472 761 -438
rect 661 -510 761 -472
rect 819 -438 919 -400
rect 819 -472 835 -438
rect 903 -472 919 -438
rect 819 -510 919 -472
rect 977 -438 1077 -400
rect 977 -472 993 -438
rect 1061 -472 1077 -438
rect 977 -510 1077 -472
rect 1135 -438 1235 -400
rect 1135 -472 1151 -438
rect 1219 -472 1235 -438
rect 1135 -510 1235 -472
rect 1293 -438 1393 -400
rect 1293 -472 1309 -438
rect 1377 -472 1393 -438
rect 1293 -510 1393 -472
rect 1451 -438 1551 -400
rect 1451 -472 1467 -438
rect 1535 -472 1551 -438
rect 1451 -510 1551 -472
rect 1609 -438 1709 -400
rect 1609 -472 1625 -438
rect 1693 -472 1709 -438
rect 1609 -510 1709 -472
rect 1767 -438 1867 -400
rect 1767 -472 1783 -438
rect 1851 -472 1867 -438
rect 1767 -510 1867 -472
rect 1925 -438 2025 -400
rect 1925 -472 1941 -438
rect 2009 -472 2025 -438
rect 1925 -510 2025 -472
rect 2083 -438 2183 -400
rect 2083 -472 2099 -438
rect 2167 -472 2183 -438
rect 2083 -510 2183 -472
rect 2241 -438 2341 -400
rect 2241 -472 2257 -438
rect 2325 -472 2341 -438
rect 2241 -510 2341 -472
rect 2399 -438 2499 -400
rect 2399 -472 2415 -438
rect 2483 -472 2499 -438
rect 2399 -510 2499 -472
rect 2557 -438 2657 -400
rect 2557 -472 2573 -438
rect 2641 -472 2657 -438
rect 2557 -510 2657 -472
rect 2715 -438 2815 -400
rect 2715 -472 2731 -438
rect 2799 -472 2815 -438
rect 2715 -510 2815 -472
rect 2873 -438 2973 -400
rect 2873 -472 2889 -438
rect 2957 -472 2973 -438
rect 2873 -510 2973 -472
rect 3031 -438 3131 -400
rect 3031 -472 3047 -438
rect 3115 -472 3131 -438
rect 3031 -510 3131 -472
rect 3189 -438 3289 -400
rect 3189 -472 3205 -438
rect 3273 -472 3289 -438
rect 3189 -510 3289 -472
rect 3347 -438 3447 -400
rect 3347 -472 3363 -438
rect 3431 -472 3447 -438
rect 3347 -510 3447 -472
rect 3505 -438 3605 -400
rect 3505 -472 3521 -438
rect 3589 -472 3605 -438
rect 3505 -510 3605 -472
rect 3663 -438 3763 -400
rect 3663 -472 3679 -438
rect 3747 -472 3763 -438
rect 3663 -510 3763 -472
rect 3821 -438 3921 -400
rect 3821 -472 3837 -438
rect 3905 -472 3921 -438
rect 3821 -510 3921 -472
rect 3979 -438 4079 -400
rect 3979 -472 3995 -438
rect 4063 -472 4079 -438
rect 3979 -510 4079 -472
rect 4137 -438 4237 -400
rect 4137 -472 4153 -438
rect 4221 -472 4237 -438
rect 4137 -510 4237 -472
rect 4295 -438 4395 -400
rect 4295 -472 4311 -438
rect 4379 -472 4395 -438
rect 4295 -510 4395 -472
rect 4453 -438 4553 -400
rect 4453 -472 4469 -438
rect 4537 -472 4553 -438
rect 4453 -510 4553 -472
rect 4611 -438 4711 -400
rect 4611 -472 4627 -438
rect 4695 -472 4711 -438
rect 4611 -510 4711 -472
rect 4769 -438 4869 -400
rect 4769 -472 4785 -438
rect 4853 -472 4869 -438
rect 4769 -510 4869 -472
rect 4927 -438 5027 -400
rect 4927 -472 4943 -438
rect 5011 -472 5027 -438
rect 4927 -510 5027 -472
rect 5085 -438 5185 -400
rect 5085 -472 5101 -438
rect 5169 -472 5185 -438
rect 5085 -510 5185 -472
rect 5243 -438 5343 -400
rect 5243 -472 5259 -438
rect 5327 -472 5343 -438
rect 5243 -510 5343 -472
rect 5401 -438 5501 -400
rect 5401 -472 5417 -438
rect 5485 -472 5501 -438
rect 5401 -510 5501 -472
rect 5559 -438 5659 -400
rect 5559 -472 5575 -438
rect 5643 -472 5659 -438
rect 5559 -510 5659 -472
rect 5717 -438 5817 -400
rect 5717 -472 5733 -438
rect 5801 -472 5817 -438
rect 5717 -510 5817 -472
rect 5875 -438 5975 -400
rect 5875 -472 5891 -438
rect 5959 -472 5975 -438
rect 5875 -510 5975 -472
rect 6033 -438 6133 -400
rect 6033 -472 6049 -438
rect 6117 -472 6133 -438
rect 6033 -510 6133 -472
rect 6191 -438 6291 -400
rect 6191 -472 6207 -438
rect 6275 -472 6291 -438
rect 6191 -510 6291 -472
rect -6291 -1348 -6191 -1310
rect -6291 -1382 -6275 -1348
rect -6207 -1382 -6191 -1348
rect -6291 -1420 -6191 -1382
rect -6133 -1348 -6033 -1310
rect -6133 -1382 -6117 -1348
rect -6049 -1382 -6033 -1348
rect -6133 -1420 -6033 -1382
rect -5975 -1348 -5875 -1310
rect -5975 -1382 -5959 -1348
rect -5891 -1382 -5875 -1348
rect -5975 -1420 -5875 -1382
rect -5817 -1348 -5717 -1310
rect -5817 -1382 -5801 -1348
rect -5733 -1382 -5717 -1348
rect -5817 -1420 -5717 -1382
rect -5659 -1348 -5559 -1310
rect -5659 -1382 -5643 -1348
rect -5575 -1382 -5559 -1348
rect -5659 -1420 -5559 -1382
rect -5501 -1348 -5401 -1310
rect -5501 -1382 -5485 -1348
rect -5417 -1382 -5401 -1348
rect -5501 -1420 -5401 -1382
rect -5343 -1348 -5243 -1310
rect -5343 -1382 -5327 -1348
rect -5259 -1382 -5243 -1348
rect -5343 -1420 -5243 -1382
rect -5185 -1348 -5085 -1310
rect -5185 -1382 -5169 -1348
rect -5101 -1382 -5085 -1348
rect -5185 -1420 -5085 -1382
rect -5027 -1348 -4927 -1310
rect -5027 -1382 -5011 -1348
rect -4943 -1382 -4927 -1348
rect -5027 -1420 -4927 -1382
rect -4869 -1348 -4769 -1310
rect -4869 -1382 -4853 -1348
rect -4785 -1382 -4769 -1348
rect -4869 -1420 -4769 -1382
rect -4711 -1348 -4611 -1310
rect -4711 -1382 -4695 -1348
rect -4627 -1382 -4611 -1348
rect -4711 -1420 -4611 -1382
rect -4553 -1348 -4453 -1310
rect -4553 -1382 -4537 -1348
rect -4469 -1382 -4453 -1348
rect -4553 -1420 -4453 -1382
rect -4395 -1348 -4295 -1310
rect -4395 -1382 -4379 -1348
rect -4311 -1382 -4295 -1348
rect -4395 -1420 -4295 -1382
rect -4237 -1348 -4137 -1310
rect -4237 -1382 -4221 -1348
rect -4153 -1382 -4137 -1348
rect -4237 -1420 -4137 -1382
rect -4079 -1348 -3979 -1310
rect -4079 -1382 -4063 -1348
rect -3995 -1382 -3979 -1348
rect -4079 -1420 -3979 -1382
rect -3921 -1348 -3821 -1310
rect -3921 -1382 -3905 -1348
rect -3837 -1382 -3821 -1348
rect -3921 -1420 -3821 -1382
rect -3763 -1348 -3663 -1310
rect -3763 -1382 -3747 -1348
rect -3679 -1382 -3663 -1348
rect -3763 -1420 -3663 -1382
rect -3605 -1348 -3505 -1310
rect -3605 -1382 -3589 -1348
rect -3521 -1382 -3505 -1348
rect -3605 -1420 -3505 -1382
rect -3447 -1348 -3347 -1310
rect -3447 -1382 -3431 -1348
rect -3363 -1382 -3347 -1348
rect -3447 -1420 -3347 -1382
rect -3289 -1348 -3189 -1310
rect -3289 -1382 -3273 -1348
rect -3205 -1382 -3189 -1348
rect -3289 -1420 -3189 -1382
rect -3131 -1348 -3031 -1310
rect -3131 -1382 -3115 -1348
rect -3047 -1382 -3031 -1348
rect -3131 -1420 -3031 -1382
rect -2973 -1348 -2873 -1310
rect -2973 -1382 -2957 -1348
rect -2889 -1382 -2873 -1348
rect -2973 -1420 -2873 -1382
rect -2815 -1348 -2715 -1310
rect -2815 -1382 -2799 -1348
rect -2731 -1382 -2715 -1348
rect -2815 -1420 -2715 -1382
rect -2657 -1348 -2557 -1310
rect -2657 -1382 -2641 -1348
rect -2573 -1382 -2557 -1348
rect -2657 -1420 -2557 -1382
rect -2499 -1348 -2399 -1310
rect -2499 -1382 -2483 -1348
rect -2415 -1382 -2399 -1348
rect -2499 -1420 -2399 -1382
rect -2341 -1348 -2241 -1310
rect -2341 -1382 -2325 -1348
rect -2257 -1382 -2241 -1348
rect -2341 -1420 -2241 -1382
rect -2183 -1348 -2083 -1310
rect -2183 -1382 -2167 -1348
rect -2099 -1382 -2083 -1348
rect -2183 -1420 -2083 -1382
rect -2025 -1348 -1925 -1310
rect -2025 -1382 -2009 -1348
rect -1941 -1382 -1925 -1348
rect -2025 -1420 -1925 -1382
rect -1867 -1348 -1767 -1310
rect -1867 -1382 -1851 -1348
rect -1783 -1382 -1767 -1348
rect -1867 -1420 -1767 -1382
rect -1709 -1348 -1609 -1310
rect -1709 -1382 -1693 -1348
rect -1625 -1382 -1609 -1348
rect -1709 -1420 -1609 -1382
rect -1551 -1348 -1451 -1310
rect -1551 -1382 -1535 -1348
rect -1467 -1382 -1451 -1348
rect -1551 -1420 -1451 -1382
rect -1393 -1348 -1293 -1310
rect -1393 -1382 -1377 -1348
rect -1309 -1382 -1293 -1348
rect -1393 -1420 -1293 -1382
rect -1235 -1348 -1135 -1310
rect -1235 -1382 -1219 -1348
rect -1151 -1382 -1135 -1348
rect -1235 -1420 -1135 -1382
rect -1077 -1348 -977 -1310
rect -1077 -1382 -1061 -1348
rect -993 -1382 -977 -1348
rect -1077 -1420 -977 -1382
rect -919 -1348 -819 -1310
rect -919 -1382 -903 -1348
rect -835 -1382 -819 -1348
rect -919 -1420 -819 -1382
rect -761 -1348 -661 -1310
rect -761 -1382 -745 -1348
rect -677 -1382 -661 -1348
rect -761 -1420 -661 -1382
rect -603 -1348 -503 -1310
rect -603 -1382 -587 -1348
rect -519 -1382 -503 -1348
rect -603 -1420 -503 -1382
rect -445 -1348 -345 -1310
rect -445 -1382 -429 -1348
rect -361 -1382 -345 -1348
rect -445 -1420 -345 -1382
rect -287 -1348 -187 -1310
rect -287 -1382 -271 -1348
rect -203 -1382 -187 -1348
rect -287 -1420 -187 -1382
rect -129 -1348 -29 -1310
rect -129 -1382 -113 -1348
rect -45 -1382 -29 -1348
rect -129 -1420 -29 -1382
rect 29 -1348 129 -1310
rect 29 -1382 45 -1348
rect 113 -1382 129 -1348
rect 29 -1420 129 -1382
rect 187 -1348 287 -1310
rect 187 -1382 203 -1348
rect 271 -1382 287 -1348
rect 187 -1420 287 -1382
rect 345 -1348 445 -1310
rect 345 -1382 361 -1348
rect 429 -1382 445 -1348
rect 345 -1420 445 -1382
rect 503 -1348 603 -1310
rect 503 -1382 519 -1348
rect 587 -1382 603 -1348
rect 503 -1420 603 -1382
rect 661 -1348 761 -1310
rect 661 -1382 677 -1348
rect 745 -1382 761 -1348
rect 661 -1420 761 -1382
rect 819 -1348 919 -1310
rect 819 -1382 835 -1348
rect 903 -1382 919 -1348
rect 819 -1420 919 -1382
rect 977 -1348 1077 -1310
rect 977 -1382 993 -1348
rect 1061 -1382 1077 -1348
rect 977 -1420 1077 -1382
rect 1135 -1348 1235 -1310
rect 1135 -1382 1151 -1348
rect 1219 -1382 1235 -1348
rect 1135 -1420 1235 -1382
rect 1293 -1348 1393 -1310
rect 1293 -1382 1309 -1348
rect 1377 -1382 1393 -1348
rect 1293 -1420 1393 -1382
rect 1451 -1348 1551 -1310
rect 1451 -1382 1467 -1348
rect 1535 -1382 1551 -1348
rect 1451 -1420 1551 -1382
rect 1609 -1348 1709 -1310
rect 1609 -1382 1625 -1348
rect 1693 -1382 1709 -1348
rect 1609 -1420 1709 -1382
rect 1767 -1348 1867 -1310
rect 1767 -1382 1783 -1348
rect 1851 -1382 1867 -1348
rect 1767 -1420 1867 -1382
rect 1925 -1348 2025 -1310
rect 1925 -1382 1941 -1348
rect 2009 -1382 2025 -1348
rect 1925 -1420 2025 -1382
rect 2083 -1348 2183 -1310
rect 2083 -1382 2099 -1348
rect 2167 -1382 2183 -1348
rect 2083 -1420 2183 -1382
rect 2241 -1348 2341 -1310
rect 2241 -1382 2257 -1348
rect 2325 -1382 2341 -1348
rect 2241 -1420 2341 -1382
rect 2399 -1348 2499 -1310
rect 2399 -1382 2415 -1348
rect 2483 -1382 2499 -1348
rect 2399 -1420 2499 -1382
rect 2557 -1348 2657 -1310
rect 2557 -1382 2573 -1348
rect 2641 -1382 2657 -1348
rect 2557 -1420 2657 -1382
rect 2715 -1348 2815 -1310
rect 2715 -1382 2731 -1348
rect 2799 -1382 2815 -1348
rect 2715 -1420 2815 -1382
rect 2873 -1348 2973 -1310
rect 2873 -1382 2889 -1348
rect 2957 -1382 2973 -1348
rect 2873 -1420 2973 -1382
rect 3031 -1348 3131 -1310
rect 3031 -1382 3047 -1348
rect 3115 -1382 3131 -1348
rect 3031 -1420 3131 -1382
rect 3189 -1348 3289 -1310
rect 3189 -1382 3205 -1348
rect 3273 -1382 3289 -1348
rect 3189 -1420 3289 -1382
rect 3347 -1348 3447 -1310
rect 3347 -1382 3363 -1348
rect 3431 -1382 3447 -1348
rect 3347 -1420 3447 -1382
rect 3505 -1348 3605 -1310
rect 3505 -1382 3521 -1348
rect 3589 -1382 3605 -1348
rect 3505 -1420 3605 -1382
rect 3663 -1348 3763 -1310
rect 3663 -1382 3679 -1348
rect 3747 -1382 3763 -1348
rect 3663 -1420 3763 -1382
rect 3821 -1348 3921 -1310
rect 3821 -1382 3837 -1348
rect 3905 -1382 3921 -1348
rect 3821 -1420 3921 -1382
rect 3979 -1348 4079 -1310
rect 3979 -1382 3995 -1348
rect 4063 -1382 4079 -1348
rect 3979 -1420 4079 -1382
rect 4137 -1348 4237 -1310
rect 4137 -1382 4153 -1348
rect 4221 -1382 4237 -1348
rect 4137 -1420 4237 -1382
rect 4295 -1348 4395 -1310
rect 4295 -1382 4311 -1348
rect 4379 -1382 4395 -1348
rect 4295 -1420 4395 -1382
rect 4453 -1348 4553 -1310
rect 4453 -1382 4469 -1348
rect 4537 -1382 4553 -1348
rect 4453 -1420 4553 -1382
rect 4611 -1348 4711 -1310
rect 4611 -1382 4627 -1348
rect 4695 -1382 4711 -1348
rect 4611 -1420 4711 -1382
rect 4769 -1348 4869 -1310
rect 4769 -1382 4785 -1348
rect 4853 -1382 4869 -1348
rect 4769 -1420 4869 -1382
rect 4927 -1348 5027 -1310
rect 4927 -1382 4943 -1348
rect 5011 -1382 5027 -1348
rect 4927 -1420 5027 -1382
rect 5085 -1348 5185 -1310
rect 5085 -1382 5101 -1348
rect 5169 -1382 5185 -1348
rect 5085 -1420 5185 -1382
rect 5243 -1348 5343 -1310
rect 5243 -1382 5259 -1348
rect 5327 -1382 5343 -1348
rect 5243 -1420 5343 -1382
rect 5401 -1348 5501 -1310
rect 5401 -1382 5417 -1348
rect 5485 -1382 5501 -1348
rect 5401 -1420 5501 -1382
rect 5559 -1348 5659 -1310
rect 5559 -1382 5575 -1348
rect 5643 -1382 5659 -1348
rect 5559 -1420 5659 -1382
rect 5717 -1348 5817 -1310
rect 5717 -1382 5733 -1348
rect 5801 -1382 5817 -1348
rect 5717 -1420 5817 -1382
rect 5875 -1348 5975 -1310
rect 5875 -1382 5891 -1348
rect 5959 -1382 5975 -1348
rect 5875 -1420 5975 -1382
rect 6033 -1348 6133 -1310
rect 6033 -1382 6049 -1348
rect 6117 -1382 6133 -1348
rect 6033 -1420 6133 -1382
rect 6191 -1348 6291 -1310
rect 6191 -1382 6207 -1348
rect 6275 -1382 6291 -1348
rect 6191 -1420 6291 -1382
rect -6291 -2258 -6191 -2220
rect -6291 -2292 -6275 -2258
rect -6207 -2292 -6191 -2258
rect -6291 -2308 -6191 -2292
rect -6133 -2258 -6033 -2220
rect -6133 -2292 -6117 -2258
rect -6049 -2292 -6033 -2258
rect -6133 -2308 -6033 -2292
rect -5975 -2258 -5875 -2220
rect -5975 -2292 -5959 -2258
rect -5891 -2292 -5875 -2258
rect -5975 -2308 -5875 -2292
rect -5817 -2258 -5717 -2220
rect -5817 -2292 -5801 -2258
rect -5733 -2292 -5717 -2258
rect -5817 -2308 -5717 -2292
rect -5659 -2258 -5559 -2220
rect -5659 -2292 -5643 -2258
rect -5575 -2292 -5559 -2258
rect -5659 -2308 -5559 -2292
rect -5501 -2258 -5401 -2220
rect -5501 -2292 -5485 -2258
rect -5417 -2292 -5401 -2258
rect -5501 -2308 -5401 -2292
rect -5343 -2258 -5243 -2220
rect -5343 -2292 -5327 -2258
rect -5259 -2292 -5243 -2258
rect -5343 -2308 -5243 -2292
rect -5185 -2258 -5085 -2220
rect -5185 -2292 -5169 -2258
rect -5101 -2292 -5085 -2258
rect -5185 -2308 -5085 -2292
rect -5027 -2258 -4927 -2220
rect -5027 -2292 -5011 -2258
rect -4943 -2292 -4927 -2258
rect -5027 -2308 -4927 -2292
rect -4869 -2258 -4769 -2220
rect -4869 -2292 -4853 -2258
rect -4785 -2292 -4769 -2258
rect -4869 -2308 -4769 -2292
rect -4711 -2258 -4611 -2220
rect -4711 -2292 -4695 -2258
rect -4627 -2292 -4611 -2258
rect -4711 -2308 -4611 -2292
rect -4553 -2258 -4453 -2220
rect -4553 -2292 -4537 -2258
rect -4469 -2292 -4453 -2258
rect -4553 -2308 -4453 -2292
rect -4395 -2258 -4295 -2220
rect -4395 -2292 -4379 -2258
rect -4311 -2292 -4295 -2258
rect -4395 -2308 -4295 -2292
rect -4237 -2258 -4137 -2220
rect -4237 -2292 -4221 -2258
rect -4153 -2292 -4137 -2258
rect -4237 -2308 -4137 -2292
rect -4079 -2258 -3979 -2220
rect -4079 -2292 -4063 -2258
rect -3995 -2292 -3979 -2258
rect -4079 -2308 -3979 -2292
rect -3921 -2258 -3821 -2220
rect -3921 -2292 -3905 -2258
rect -3837 -2292 -3821 -2258
rect -3921 -2308 -3821 -2292
rect -3763 -2258 -3663 -2220
rect -3763 -2292 -3747 -2258
rect -3679 -2292 -3663 -2258
rect -3763 -2308 -3663 -2292
rect -3605 -2258 -3505 -2220
rect -3605 -2292 -3589 -2258
rect -3521 -2292 -3505 -2258
rect -3605 -2308 -3505 -2292
rect -3447 -2258 -3347 -2220
rect -3447 -2292 -3431 -2258
rect -3363 -2292 -3347 -2258
rect -3447 -2308 -3347 -2292
rect -3289 -2258 -3189 -2220
rect -3289 -2292 -3273 -2258
rect -3205 -2292 -3189 -2258
rect -3289 -2308 -3189 -2292
rect -3131 -2258 -3031 -2220
rect -3131 -2292 -3115 -2258
rect -3047 -2292 -3031 -2258
rect -3131 -2308 -3031 -2292
rect -2973 -2258 -2873 -2220
rect -2973 -2292 -2957 -2258
rect -2889 -2292 -2873 -2258
rect -2973 -2308 -2873 -2292
rect -2815 -2258 -2715 -2220
rect -2815 -2292 -2799 -2258
rect -2731 -2292 -2715 -2258
rect -2815 -2308 -2715 -2292
rect -2657 -2258 -2557 -2220
rect -2657 -2292 -2641 -2258
rect -2573 -2292 -2557 -2258
rect -2657 -2308 -2557 -2292
rect -2499 -2258 -2399 -2220
rect -2499 -2292 -2483 -2258
rect -2415 -2292 -2399 -2258
rect -2499 -2308 -2399 -2292
rect -2341 -2258 -2241 -2220
rect -2341 -2292 -2325 -2258
rect -2257 -2292 -2241 -2258
rect -2341 -2308 -2241 -2292
rect -2183 -2258 -2083 -2220
rect -2183 -2292 -2167 -2258
rect -2099 -2292 -2083 -2258
rect -2183 -2308 -2083 -2292
rect -2025 -2258 -1925 -2220
rect -2025 -2292 -2009 -2258
rect -1941 -2292 -1925 -2258
rect -2025 -2308 -1925 -2292
rect -1867 -2258 -1767 -2220
rect -1867 -2292 -1851 -2258
rect -1783 -2292 -1767 -2258
rect -1867 -2308 -1767 -2292
rect -1709 -2258 -1609 -2220
rect -1709 -2292 -1693 -2258
rect -1625 -2292 -1609 -2258
rect -1709 -2308 -1609 -2292
rect -1551 -2258 -1451 -2220
rect -1551 -2292 -1535 -2258
rect -1467 -2292 -1451 -2258
rect -1551 -2308 -1451 -2292
rect -1393 -2258 -1293 -2220
rect -1393 -2292 -1377 -2258
rect -1309 -2292 -1293 -2258
rect -1393 -2308 -1293 -2292
rect -1235 -2258 -1135 -2220
rect -1235 -2292 -1219 -2258
rect -1151 -2292 -1135 -2258
rect -1235 -2308 -1135 -2292
rect -1077 -2258 -977 -2220
rect -1077 -2292 -1061 -2258
rect -993 -2292 -977 -2258
rect -1077 -2308 -977 -2292
rect -919 -2258 -819 -2220
rect -919 -2292 -903 -2258
rect -835 -2292 -819 -2258
rect -919 -2308 -819 -2292
rect -761 -2258 -661 -2220
rect -761 -2292 -745 -2258
rect -677 -2292 -661 -2258
rect -761 -2308 -661 -2292
rect -603 -2258 -503 -2220
rect -603 -2292 -587 -2258
rect -519 -2292 -503 -2258
rect -603 -2308 -503 -2292
rect -445 -2258 -345 -2220
rect -445 -2292 -429 -2258
rect -361 -2292 -345 -2258
rect -445 -2308 -345 -2292
rect -287 -2258 -187 -2220
rect -287 -2292 -271 -2258
rect -203 -2292 -187 -2258
rect -287 -2308 -187 -2292
rect -129 -2258 -29 -2220
rect -129 -2292 -113 -2258
rect -45 -2292 -29 -2258
rect -129 -2308 -29 -2292
rect 29 -2258 129 -2220
rect 29 -2292 45 -2258
rect 113 -2292 129 -2258
rect 29 -2308 129 -2292
rect 187 -2258 287 -2220
rect 187 -2292 203 -2258
rect 271 -2292 287 -2258
rect 187 -2308 287 -2292
rect 345 -2258 445 -2220
rect 345 -2292 361 -2258
rect 429 -2292 445 -2258
rect 345 -2308 445 -2292
rect 503 -2258 603 -2220
rect 503 -2292 519 -2258
rect 587 -2292 603 -2258
rect 503 -2308 603 -2292
rect 661 -2258 761 -2220
rect 661 -2292 677 -2258
rect 745 -2292 761 -2258
rect 661 -2308 761 -2292
rect 819 -2258 919 -2220
rect 819 -2292 835 -2258
rect 903 -2292 919 -2258
rect 819 -2308 919 -2292
rect 977 -2258 1077 -2220
rect 977 -2292 993 -2258
rect 1061 -2292 1077 -2258
rect 977 -2308 1077 -2292
rect 1135 -2258 1235 -2220
rect 1135 -2292 1151 -2258
rect 1219 -2292 1235 -2258
rect 1135 -2308 1235 -2292
rect 1293 -2258 1393 -2220
rect 1293 -2292 1309 -2258
rect 1377 -2292 1393 -2258
rect 1293 -2308 1393 -2292
rect 1451 -2258 1551 -2220
rect 1451 -2292 1467 -2258
rect 1535 -2292 1551 -2258
rect 1451 -2308 1551 -2292
rect 1609 -2258 1709 -2220
rect 1609 -2292 1625 -2258
rect 1693 -2292 1709 -2258
rect 1609 -2308 1709 -2292
rect 1767 -2258 1867 -2220
rect 1767 -2292 1783 -2258
rect 1851 -2292 1867 -2258
rect 1767 -2308 1867 -2292
rect 1925 -2258 2025 -2220
rect 1925 -2292 1941 -2258
rect 2009 -2292 2025 -2258
rect 1925 -2308 2025 -2292
rect 2083 -2258 2183 -2220
rect 2083 -2292 2099 -2258
rect 2167 -2292 2183 -2258
rect 2083 -2308 2183 -2292
rect 2241 -2258 2341 -2220
rect 2241 -2292 2257 -2258
rect 2325 -2292 2341 -2258
rect 2241 -2308 2341 -2292
rect 2399 -2258 2499 -2220
rect 2399 -2292 2415 -2258
rect 2483 -2292 2499 -2258
rect 2399 -2308 2499 -2292
rect 2557 -2258 2657 -2220
rect 2557 -2292 2573 -2258
rect 2641 -2292 2657 -2258
rect 2557 -2308 2657 -2292
rect 2715 -2258 2815 -2220
rect 2715 -2292 2731 -2258
rect 2799 -2292 2815 -2258
rect 2715 -2308 2815 -2292
rect 2873 -2258 2973 -2220
rect 2873 -2292 2889 -2258
rect 2957 -2292 2973 -2258
rect 2873 -2308 2973 -2292
rect 3031 -2258 3131 -2220
rect 3031 -2292 3047 -2258
rect 3115 -2292 3131 -2258
rect 3031 -2308 3131 -2292
rect 3189 -2258 3289 -2220
rect 3189 -2292 3205 -2258
rect 3273 -2292 3289 -2258
rect 3189 -2308 3289 -2292
rect 3347 -2258 3447 -2220
rect 3347 -2292 3363 -2258
rect 3431 -2292 3447 -2258
rect 3347 -2308 3447 -2292
rect 3505 -2258 3605 -2220
rect 3505 -2292 3521 -2258
rect 3589 -2292 3605 -2258
rect 3505 -2308 3605 -2292
rect 3663 -2258 3763 -2220
rect 3663 -2292 3679 -2258
rect 3747 -2292 3763 -2258
rect 3663 -2308 3763 -2292
rect 3821 -2258 3921 -2220
rect 3821 -2292 3837 -2258
rect 3905 -2292 3921 -2258
rect 3821 -2308 3921 -2292
rect 3979 -2258 4079 -2220
rect 3979 -2292 3995 -2258
rect 4063 -2292 4079 -2258
rect 3979 -2308 4079 -2292
rect 4137 -2258 4237 -2220
rect 4137 -2292 4153 -2258
rect 4221 -2292 4237 -2258
rect 4137 -2308 4237 -2292
rect 4295 -2258 4395 -2220
rect 4295 -2292 4311 -2258
rect 4379 -2292 4395 -2258
rect 4295 -2308 4395 -2292
rect 4453 -2258 4553 -2220
rect 4453 -2292 4469 -2258
rect 4537 -2292 4553 -2258
rect 4453 -2308 4553 -2292
rect 4611 -2258 4711 -2220
rect 4611 -2292 4627 -2258
rect 4695 -2292 4711 -2258
rect 4611 -2308 4711 -2292
rect 4769 -2258 4869 -2220
rect 4769 -2292 4785 -2258
rect 4853 -2292 4869 -2258
rect 4769 -2308 4869 -2292
rect 4927 -2258 5027 -2220
rect 4927 -2292 4943 -2258
rect 5011 -2292 5027 -2258
rect 4927 -2308 5027 -2292
rect 5085 -2258 5185 -2220
rect 5085 -2292 5101 -2258
rect 5169 -2292 5185 -2258
rect 5085 -2308 5185 -2292
rect 5243 -2258 5343 -2220
rect 5243 -2292 5259 -2258
rect 5327 -2292 5343 -2258
rect 5243 -2308 5343 -2292
rect 5401 -2258 5501 -2220
rect 5401 -2292 5417 -2258
rect 5485 -2292 5501 -2258
rect 5401 -2308 5501 -2292
rect 5559 -2258 5659 -2220
rect 5559 -2292 5575 -2258
rect 5643 -2292 5659 -2258
rect 5559 -2308 5659 -2292
rect 5717 -2258 5817 -2220
rect 5717 -2292 5733 -2258
rect 5801 -2292 5817 -2258
rect 5717 -2308 5817 -2292
rect 5875 -2258 5975 -2220
rect 5875 -2292 5891 -2258
rect 5959 -2292 5975 -2258
rect 5875 -2308 5975 -2292
rect 6033 -2258 6133 -2220
rect 6033 -2292 6049 -2258
rect 6117 -2292 6133 -2258
rect 6033 -2308 6133 -2292
rect 6191 -2258 6291 -2220
rect 6191 -2292 6207 -2258
rect 6275 -2292 6291 -2258
rect 6191 -2308 6291 -2292
<< polycont >>
rect -6275 2258 -6207 2292
rect -6117 2258 -6049 2292
rect -5959 2258 -5891 2292
rect -5801 2258 -5733 2292
rect -5643 2258 -5575 2292
rect -5485 2258 -5417 2292
rect -5327 2258 -5259 2292
rect -5169 2258 -5101 2292
rect -5011 2258 -4943 2292
rect -4853 2258 -4785 2292
rect -4695 2258 -4627 2292
rect -4537 2258 -4469 2292
rect -4379 2258 -4311 2292
rect -4221 2258 -4153 2292
rect -4063 2258 -3995 2292
rect -3905 2258 -3837 2292
rect -3747 2258 -3679 2292
rect -3589 2258 -3521 2292
rect -3431 2258 -3363 2292
rect -3273 2258 -3205 2292
rect -3115 2258 -3047 2292
rect -2957 2258 -2889 2292
rect -2799 2258 -2731 2292
rect -2641 2258 -2573 2292
rect -2483 2258 -2415 2292
rect -2325 2258 -2257 2292
rect -2167 2258 -2099 2292
rect -2009 2258 -1941 2292
rect -1851 2258 -1783 2292
rect -1693 2258 -1625 2292
rect -1535 2258 -1467 2292
rect -1377 2258 -1309 2292
rect -1219 2258 -1151 2292
rect -1061 2258 -993 2292
rect -903 2258 -835 2292
rect -745 2258 -677 2292
rect -587 2258 -519 2292
rect -429 2258 -361 2292
rect -271 2258 -203 2292
rect -113 2258 -45 2292
rect 45 2258 113 2292
rect 203 2258 271 2292
rect 361 2258 429 2292
rect 519 2258 587 2292
rect 677 2258 745 2292
rect 835 2258 903 2292
rect 993 2258 1061 2292
rect 1151 2258 1219 2292
rect 1309 2258 1377 2292
rect 1467 2258 1535 2292
rect 1625 2258 1693 2292
rect 1783 2258 1851 2292
rect 1941 2258 2009 2292
rect 2099 2258 2167 2292
rect 2257 2258 2325 2292
rect 2415 2258 2483 2292
rect 2573 2258 2641 2292
rect 2731 2258 2799 2292
rect 2889 2258 2957 2292
rect 3047 2258 3115 2292
rect 3205 2258 3273 2292
rect 3363 2258 3431 2292
rect 3521 2258 3589 2292
rect 3679 2258 3747 2292
rect 3837 2258 3905 2292
rect 3995 2258 4063 2292
rect 4153 2258 4221 2292
rect 4311 2258 4379 2292
rect 4469 2258 4537 2292
rect 4627 2258 4695 2292
rect 4785 2258 4853 2292
rect 4943 2258 5011 2292
rect 5101 2258 5169 2292
rect 5259 2258 5327 2292
rect 5417 2258 5485 2292
rect 5575 2258 5643 2292
rect 5733 2258 5801 2292
rect 5891 2258 5959 2292
rect 6049 2258 6117 2292
rect 6207 2258 6275 2292
rect -6275 1348 -6207 1382
rect -6117 1348 -6049 1382
rect -5959 1348 -5891 1382
rect -5801 1348 -5733 1382
rect -5643 1348 -5575 1382
rect -5485 1348 -5417 1382
rect -5327 1348 -5259 1382
rect -5169 1348 -5101 1382
rect -5011 1348 -4943 1382
rect -4853 1348 -4785 1382
rect -4695 1348 -4627 1382
rect -4537 1348 -4469 1382
rect -4379 1348 -4311 1382
rect -4221 1348 -4153 1382
rect -4063 1348 -3995 1382
rect -3905 1348 -3837 1382
rect -3747 1348 -3679 1382
rect -3589 1348 -3521 1382
rect -3431 1348 -3363 1382
rect -3273 1348 -3205 1382
rect -3115 1348 -3047 1382
rect -2957 1348 -2889 1382
rect -2799 1348 -2731 1382
rect -2641 1348 -2573 1382
rect -2483 1348 -2415 1382
rect -2325 1348 -2257 1382
rect -2167 1348 -2099 1382
rect -2009 1348 -1941 1382
rect -1851 1348 -1783 1382
rect -1693 1348 -1625 1382
rect -1535 1348 -1467 1382
rect -1377 1348 -1309 1382
rect -1219 1348 -1151 1382
rect -1061 1348 -993 1382
rect -903 1348 -835 1382
rect -745 1348 -677 1382
rect -587 1348 -519 1382
rect -429 1348 -361 1382
rect -271 1348 -203 1382
rect -113 1348 -45 1382
rect 45 1348 113 1382
rect 203 1348 271 1382
rect 361 1348 429 1382
rect 519 1348 587 1382
rect 677 1348 745 1382
rect 835 1348 903 1382
rect 993 1348 1061 1382
rect 1151 1348 1219 1382
rect 1309 1348 1377 1382
rect 1467 1348 1535 1382
rect 1625 1348 1693 1382
rect 1783 1348 1851 1382
rect 1941 1348 2009 1382
rect 2099 1348 2167 1382
rect 2257 1348 2325 1382
rect 2415 1348 2483 1382
rect 2573 1348 2641 1382
rect 2731 1348 2799 1382
rect 2889 1348 2957 1382
rect 3047 1348 3115 1382
rect 3205 1348 3273 1382
rect 3363 1348 3431 1382
rect 3521 1348 3589 1382
rect 3679 1348 3747 1382
rect 3837 1348 3905 1382
rect 3995 1348 4063 1382
rect 4153 1348 4221 1382
rect 4311 1348 4379 1382
rect 4469 1348 4537 1382
rect 4627 1348 4695 1382
rect 4785 1348 4853 1382
rect 4943 1348 5011 1382
rect 5101 1348 5169 1382
rect 5259 1348 5327 1382
rect 5417 1348 5485 1382
rect 5575 1348 5643 1382
rect 5733 1348 5801 1382
rect 5891 1348 5959 1382
rect 6049 1348 6117 1382
rect 6207 1348 6275 1382
rect -6275 438 -6207 472
rect -6117 438 -6049 472
rect -5959 438 -5891 472
rect -5801 438 -5733 472
rect -5643 438 -5575 472
rect -5485 438 -5417 472
rect -5327 438 -5259 472
rect -5169 438 -5101 472
rect -5011 438 -4943 472
rect -4853 438 -4785 472
rect -4695 438 -4627 472
rect -4537 438 -4469 472
rect -4379 438 -4311 472
rect -4221 438 -4153 472
rect -4063 438 -3995 472
rect -3905 438 -3837 472
rect -3747 438 -3679 472
rect -3589 438 -3521 472
rect -3431 438 -3363 472
rect -3273 438 -3205 472
rect -3115 438 -3047 472
rect -2957 438 -2889 472
rect -2799 438 -2731 472
rect -2641 438 -2573 472
rect -2483 438 -2415 472
rect -2325 438 -2257 472
rect -2167 438 -2099 472
rect -2009 438 -1941 472
rect -1851 438 -1783 472
rect -1693 438 -1625 472
rect -1535 438 -1467 472
rect -1377 438 -1309 472
rect -1219 438 -1151 472
rect -1061 438 -993 472
rect -903 438 -835 472
rect -745 438 -677 472
rect -587 438 -519 472
rect -429 438 -361 472
rect -271 438 -203 472
rect -113 438 -45 472
rect 45 438 113 472
rect 203 438 271 472
rect 361 438 429 472
rect 519 438 587 472
rect 677 438 745 472
rect 835 438 903 472
rect 993 438 1061 472
rect 1151 438 1219 472
rect 1309 438 1377 472
rect 1467 438 1535 472
rect 1625 438 1693 472
rect 1783 438 1851 472
rect 1941 438 2009 472
rect 2099 438 2167 472
rect 2257 438 2325 472
rect 2415 438 2483 472
rect 2573 438 2641 472
rect 2731 438 2799 472
rect 2889 438 2957 472
rect 3047 438 3115 472
rect 3205 438 3273 472
rect 3363 438 3431 472
rect 3521 438 3589 472
rect 3679 438 3747 472
rect 3837 438 3905 472
rect 3995 438 4063 472
rect 4153 438 4221 472
rect 4311 438 4379 472
rect 4469 438 4537 472
rect 4627 438 4695 472
rect 4785 438 4853 472
rect 4943 438 5011 472
rect 5101 438 5169 472
rect 5259 438 5327 472
rect 5417 438 5485 472
rect 5575 438 5643 472
rect 5733 438 5801 472
rect 5891 438 5959 472
rect 6049 438 6117 472
rect 6207 438 6275 472
rect -6275 -472 -6207 -438
rect -6117 -472 -6049 -438
rect -5959 -472 -5891 -438
rect -5801 -472 -5733 -438
rect -5643 -472 -5575 -438
rect -5485 -472 -5417 -438
rect -5327 -472 -5259 -438
rect -5169 -472 -5101 -438
rect -5011 -472 -4943 -438
rect -4853 -472 -4785 -438
rect -4695 -472 -4627 -438
rect -4537 -472 -4469 -438
rect -4379 -472 -4311 -438
rect -4221 -472 -4153 -438
rect -4063 -472 -3995 -438
rect -3905 -472 -3837 -438
rect -3747 -472 -3679 -438
rect -3589 -472 -3521 -438
rect -3431 -472 -3363 -438
rect -3273 -472 -3205 -438
rect -3115 -472 -3047 -438
rect -2957 -472 -2889 -438
rect -2799 -472 -2731 -438
rect -2641 -472 -2573 -438
rect -2483 -472 -2415 -438
rect -2325 -472 -2257 -438
rect -2167 -472 -2099 -438
rect -2009 -472 -1941 -438
rect -1851 -472 -1783 -438
rect -1693 -472 -1625 -438
rect -1535 -472 -1467 -438
rect -1377 -472 -1309 -438
rect -1219 -472 -1151 -438
rect -1061 -472 -993 -438
rect -903 -472 -835 -438
rect -745 -472 -677 -438
rect -587 -472 -519 -438
rect -429 -472 -361 -438
rect -271 -472 -203 -438
rect -113 -472 -45 -438
rect 45 -472 113 -438
rect 203 -472 271 -438
rect 361 -472 429 -438
rect 519 -472 587 -438
rect 677 -472 745 -438
rect 835 -472 903 -438
rect 993 -472 1061 -438
rect 1151 -472 1219 -438
rect 1309 -472 1377 -438
rect 1467 -472 1535 -438
rect 1625 -472 1693 -438
rect 1783 -472 1851 -438
rect 1941 -472 2009 -438
rect 2099 -472 2167 -438
rect 2257 -472 2325 -438
rect 2415 -472 2483 -438
rect 2573 -472 2641 -438
rect 2731 -472 2799 -438
rect 2889 -472 2957 -438
rect 3047 -472 3115 -438
rect 3205 -472 3273 -438
rect 3363 -472 3431 -438
rect 3521 -472 3589 -438
rect 3679 -472 3747 -438
rect 3837 -472 3905 -438
rect 3995 -472 4063 -438
rect 4153 -472 4221 -438
rect 4311 -472 4379 -438
rect 4469 -472 4537 -438
rect 4627 -472 4695 -438
rect 4785 -472 4853 -438
rect 4943 -472 5011 -438
rect 5101 -472 5169 -438
rect 5259 -472 5327 -438
rect 5417 -472 5485 -438
rect 5575 -472 5643 -438
rect 5733 -472 5801 -438
rect 5891 -472 5959 -438
rect 6049 -472 6117 -438
rect 6207 -472 6275 -438
rect -6275 -1382 -6207 -1348
rect -6117 -1382 -6049 -1348
rect -5959 -1382 -5891 -1348
rect -5801 -1382 -5733 -1348
rect -5643 -1382 -5575 -1348
rect -5485 -1382 -5417 -1348
rect -5327 -1382 -5259 -1348
rect -5169 -1382 -5101 -1348
rect -5011 -1382 -4943 -1348
rect -4853 -1382 -4785 -1348
rect -4695 -1382 -4627 -1348
rect -4537 -1382 -4469 -1348
rect -4379 -1382 -4311 -1348
rect -4221 -1382 -4153 -1348
rect -4063 -1382 -3995 -1348
rect -3905 -1382 -3837 -1348
rect -3747 -1382 -3679 -1348
rect -3589 -1382 -3521 -1348
rect -3431 -1382 -3363 -1348
rect -3273 -1382 -3205 -1348
rect -3115 -1382 -3047 -1348
rect -2957 -1382 -2889 -1348
rect -2799 -1382 -2731 -1348
rect -2641 -1382 -2573 -1348
rect -2483 -1382 -2415 -1348
rect -2325 -1382 -2257 -1348
rect -2167 -1382 -2099 -1348
rect -2009 -1382 -1941 -1348
rect -1851 -1382 -1783 -1348
rect -1693 -1382 -1625 -1348
rect -1535 -1382 -1467 -1348
rect -1377 -1382 -1309 -1348
rect -1219 -1382 -1151 -1348
rect -1061 -1382 -993 -1348
rect -903 -1382 -835 -1348
rect -745 -1382 -677 -1348
rect -587 -1382 -519 -1348
rect -429 -1382 -361 -1348
rect -271 -1382 -203 -1348
rect -113 -1382 -45 -1348
rect 45 -1382 113 -1348
rect 203 -1382 271 -1348
rect 361 -1382 429 -1348
rect 519 -1382 587 -1348
rect 677 -1382 745 -1348
rect 835 -1382 903 -1348
rect 993 -1382 1061 -1348
rect 1151 -1382 1219 -1348
rect 1309 -1382 1377 -1348
rect 1467 -1382 1535 -1348
rect 1625 -1382 1693 -1348
rect 1783 -1382 1851 -1348
rect 1941 -1382 2009 -1348
rect 2099 -1382 2167 -1348
rect 2257 -1382 2325 -1348
rect 2415 -1382 2483 -1348
rect 2573 -1382 2641 -1348
rect 2731 -1382 2799 -1348
rect 2889 -1382 2957 -1348
rect 3047 -1382 3115 -1348
rect 3205 -1382 3273 -1348
rect 3363 -1382 3431 -1348
rect 3521 -1382 3589 -1348
rect 3679 -1382 3747 -1348
rect 3837 -1382 3905 -1348
rect 3995 -1382 4063 -1348
rect 4153 -1382 4221 -1348
rect 4311 -1382 4379 -1348
rect 4469 -1382 4537 -1348
rect 4627 -1382 4695 -1348
rect 4785 -1382 4853 -1348
rect 4943 -1382 5011 -1348
rect 5101 -1382 5169 -1348
rect 5259 -1382 5327 -1348
rect 5417 -1382 5485 -1348
rect 5575 -1382 5643 -1348
rect 5733 -1382 5801 -1348
rect 5891 -1382 5959 -1348
rect 6049 -1382 6117 -1348
rect 6207 -1382 6275 -1348
rect -6275 -2292 -6207 -2258
rect -6117 -2292 -6049 -2258
rect -5959 -2292 -5891 -2258
rect -5801 -2292 -5733 -2258
rect -5643 -2292 -5575 -2258
rect -5485 -2292 -5417 -2258
rect -5327 -2292 -5259 -2258
rect -5169 -2292 -5101 -2258
rect -5011 -2292 -4943 -2258
rect -4853 -2292 -4785 -2258
rect -4695 -2292 -4627 -2258
rect -4537 -2292 -4469 -2258
rect -4379 -2292 -4311 -2258
rect -4221 -2292 -4153 -2258
rect -4063 -2292 -3995 -2258
rect -3905 -2292 -3837 -2258
rect -3747 -2292 -3679 -2258
rect -3589 -2292 -3521 -2258
rect -3431 -2292 -3363 -2258
rect -3273 -2292 -3205 -2258
rect -3115 -2292 -3047 -2258
rect -2957 -2292 -2889 -2258
rect -2799 -2292 -2731 -2258
rect -2641 -2292 -2573 -2258
rect -2483 -2292 -2415 -2258
rect -2325 -2292 -2257 -2258
rect -2167 -2292 -2099 -2258
rect -2009 -2292 -1941 -2258
rect -1851 -2292 -1783 -2258
rect -1693 -2292 -1625 -2258
rect -1535 -2292 -1467 -2258
rect -1377 -2292 -1309 -2258
rect -1219 -2292 -1151 -2258
rect -1061 -2292 -993 -2258
rect -903 -2292 -835 -2258
rect -745 -2292 -677 -2258
rect -587 -2292 -519 -2258
rect -429 -2292 -361 -2258
rect -271 -2292 -203 -2258
rect -113 -2292 -45 -2258
rect 45 -2292 113 -2258
rect 203 -2292 271 -2258
rect 361 -2292 429 -2258
rect 519 -2292 587 -2258
rect 677 -2292 745 -2258
rect 835 -2292 903 -2258
rect 993 -2292 1061 -2258
rect 1151 -2292 1219 -2258
rect 1309 -2292 1377 -2258
rect 1467 -2292 1535 -2258
rect 1625 -2292 1693 -2258
rect 1783 -2292 1851 -2258
rect 1941 -2292 2009 -2258
rect 2099 -2292 2167 -2258
rect 2257 -2292 2325 -2258
rect 2415 -2292 2483 -2258
rect 2573 -2292 2641 -2258
rect 2731 -2292 2799 -2258
rect 2889 -2292 2957 -2258
rect 3047 -2292 3115 -2258
rect 3205 -2292 3273 -2258
rect 3363 -2292 3431 -2258
rect 3521 -2292 3589 -2258
rect 3679 -2292 3747 -2258
rect 3837 -2292 3905 -2258
rect 3995 -2292 4063 -2258
rect 4153 -2292 4221 -2258
rect 4311 -2292 4379 -2258
rect 4469 -2292 4537 -2258
rect 4627 -2292 4695 -2258
rect 4785 -2292 4853 -2258
rect 4943 -2292 5011 -2258
rect 5101 -2292 5169 -2258
rect 5259 -2292 5327 -2258
rect 5417 -2292 5485 -2258
rect 5575 -2292 5643 -2258
rect 5733 -2292 5801 -2258
rect 5891 -2292 5959 -2258
rect 6049 -2292 6117 -2258
rect 6207 -2292 6275 -2258
<< locali >>
rect -6471 2396 -6375 2430
rect 6375 2396 6471 2430
rect -6471 2334 -6437 2396
rect 6437 2334 6471 2396
rect -6291 2258 -6275 2292
rect -6207 2258 -6191 2292
rect -6133 2258 -6117 2292
rect -6049 2258 -6033 2292
rect -5975 2258 -5959 2292
rect -5891 2258 -5875 2292
rect -5817 2258 -5801 2292
rect -5733 2258 -5717 2292
rect -5659 2258 -5643 2292
rect -5575 2258 -5559 2292
rect -5501 2258 -5485 2292
rect -5417 2258 -5401 2292
rect -5343 2258 -5327 2292
rect -5259 2258 -5243 2292
rect -5185 2258 -5169 2292
rect -5101 2258 -5085 2292
rect -5027 2258 -5011 2292
rect -4943 2258 -4927 2292
rect -4869 2258 -4853 2292
rect -4785 2258 -4769 2292
rect -4711 2258 -4695 2292
rect -4627 2258 -4611 2292
rect -4553 2258 -4537 2292
rect -4469 2258 -4453 2292
rect -4395 2258 -4379 2292
rect -4311 2258 -4295 2292
rect -4237 2258 -4221 2292
rect -4153 2258 -4137 2292
rect -4079 2258 -4063 2292
rect -3995 2258 -3979 2292
rect -3921 2258 -3905 2292
rect -3837 2258 -3821 2292
rect -3763 2258 -3747 2292
rect -3679 2258 -3663 2292
rect -3605 2258 -3589 2292
rect -3521 2258 -3505 2292
rect -3447 2258 -3431 2292
rect -3363 2258 -3347 2292
rect -3289 2258 -3273 2292
rect -3205 2258 -3189 2292
rect -3131 2258 -3115 2292
rect -3047 2258 -3031 2292
rect -2973 2258 -2957 2292
rect -2889 2258 -2873 2292
rect -2815 2258 -2799 2292
rect -2731 2258 -2715 2292
rect -2657 2258 -2641 2292
rect -2573 2258 -2557 2292
rect -2499 2258 -2483 2292
rect -2415 2258 -2399 2292
rect -2341 2258 -2325 2292
rect -2257 2258 -2241 2292
rect -2183 2258 -2167 2292
rect -2099 2258 -2083 2292
rect -2025 2258 -2009 2292
rect -1941 2258 -1925 2292
rect -1867 2258 -1851 2292
rect -1783 2258 -1767 2292
rect -1709 2258 -1693 2292
rect -1625 2258 -1609 2292
rect -1551 2258 -1535 2292
rect -1467 2258 -1451 2292
rect -1393 2258 -1377 2292
rect -1309 2258 -1293 2292
rect -1235 2258 -1219 2292
rect -1151 2258 -1135 2292
rect -1077 2258 -1061 2292
rect -993 2258 -977 2292
rect -919 2258 -903 2292
rect -835 2258 -819 2292
rect -761 2258 -745 2292
rect -677 2258 -661 2292
rect -603 2258 -587 2292
rect -519 2258 -503 2292
rect -445 2258 -429 2292
rect -361 2258 -345 2292
rect -287 2258 -271 2292
rect -203 2258 -187 2292
rect -129 2258 -113 2292
rect -45 2258 -29 2292
rect 29 2258 45 2292
rect 113 2258 129 2292
rect 187 2258 203 2292
rect 271 2258 287 2292
rect 345 2258 361 2292
rect 429 2258 445 2292
rect 503 2258 519 2292
rect 587 2258 603 2292
rect 661 2258 677 2292
rect 745 2258 761 2292
rect 819 2258 835 2292
rect 903 2258 919 2292
rect 977 2258 993 2292
rect 1061 2258 1077 2292
rect 1135 2258 1151 2292
rect 1219 2258 1235 2292
rect 1293 2258 1309 2292
rect 1377 2258 1393 2292
rect 1451 2258 1467 2292
rect 1535 2258 1551 2292
rect 1609 2258 1625 2292
rect 1693 2258 1709 2292
rect 1767 2258 1783 2292
rect 1851 2258 1867 2292
rect 1925 2258 1941 2292
rect 2009 2258 2025 2292
rect 2083 2258 2099 2292
rect 2167 2258 2183 2292
rect 2241 2258 2257 2292
rect 2325 2258 2341 2292
rect 2399 2258 2415 2292
rect 2483 2258 2499 2292
rect 2557 2258 2573 2292
rect 2641 2258 2657 2292
rect 2715 2258 2731 2292
rect 2799 2258 2815 2292
rect 2873 2258 2889 2292
rect 2957 2258 2973 2292
rect 3031 2258 3047 2292
rect 3115 2258 3131 2292
rect 3189 2258 3205 2292
rect 3273 2258 3289 2292
rect 3347 2258 3363 2292
rect 3431 2258 3447 2292
rect 3505 2258 3521 2292
rect 3589 2258 3605 2292
rect 3663 2258 3679 2292
rect 3747 2258 3763 2292
rect 3821 2258 3837 2292
rect 3905 2258 3921 2292
rect 3979 2258 3995 2292
rect 4063 2258 4079 2292
rect 4137 2258 4153 2292
rect 4221 2258 4237 2292
rect 4295 2258 4311 2292
rect 4379 2258 4395 2292
rect 4453 2258 4469 2292
rect 4537 2258 4553 2292
rect 4611 2258 4627 2292
rect 4695 2258 4711 2292
rect 4769 2258 4785 2292
rect 4853 2258 4869 2292
rect 4927 2258 4943 2292
rect 5011 2258 5027 2292
rect 5085 2258 5101 2292
rect 5169 2258 5185 2292
rect 5243 2258 5259 2292
rect 5327 2258 5343 2292
rect 5401 2258 5417 2292
rect 5485 2258 5501 2292
rect 5559 2258 5575 2292
rect 5643 2258 5659 2292
rect 5717 2258 5733 2292
rect 5801 2258 5817 2292
rect 5875 2258 5891 2292
rect 5959 2258 5975 2292
rect 6033 2258 6049 2292
rect 6117 2258 6133 2292
rect 6191 2258 6207 2292
rect 6275 2258 6291 2292
rect -6337 2208 -6303 2224
rect -6337 1416 -6303 1432
rect -6179 2208 -6145 2224
rect -6179 1416 -6145 1432
rect -6021 2208 -5987 2224
rect -6021 1416 -5987 1432
rect -5863 2208 -5829 2224
rect -5863 1416 -5829 1432
rect -5705 2208 -5671 2224
rect -5705 1416 -5671 1432
rect -5547 2208 -5513 2224
rect -5547 1416 -5513 1432
rect -5389 2208 -5355 2224
rect -5389 1416 -5355 1432
rect -5231 2208 -5197 2224
rect -5231 1416 -5197 1432
rect -5073 2208 -5039 2224
rect -5073 1416 -5039 1432
rect -4915 2208 -4881 2224
rect -4915 1416 -4881 1432
rect -4757 2208 -4723 2224
rect -4757 1416 -4723 1432
rect -4599 2208 -4565 2224
rect -4599 1416 -4565 1432
rect -4441 2208 -4407 2224
rect -4441 1416 -4407 1432
rect -4283 2208 -4249 2224
rect -4283 1416 -4249 1432
rect -4125 2208 -4091 2224
rect -4125 1416 -4091 1432
rect -3967 2208 -3933 2224
rect -3967 1416 -3933 1432
rect -3809 2208 -3775 2224
rect -3809 1416 -3775 1432
rect -3651 2208 -3617 2224
rect -3651 1416 -3617 1432
rect -3493 2208 -3459 2224
rect -3493 1416 -3459 1432
rect -3335 2208 -3301 2224
rect -3335 1416 -3301 1432
rect -3177 2208 -3143 2224
rect -3177 1416 -3143 1432
rect -3019 2208 -2985 2224
rect -3019 1416 -2985 1432
rect -2861 2208 -2827 2224
rect -2861 1416 -2827 1432
rect -2703 2208 -2669 2224
rect -2703 1416 -2669 1432
rect -2545 2208 -2511 2224
rect -2545 1416 -2511 1432
rect -2387 2208 -2353 2224
rect -2387 1416 -2353 1432
rect -2229 2208 -2195 2224
rect -2229 1416 -2195 1432
rect -2071 2208 -2037 2224
rect -2071 1416 -2037 1432
rect -1913 2208 -1879 2224
rect -1913 1416 -1879 1432
rect -1755 2208 -1721 2224
rect -1755 1416 -1721 1432
rect -1597 2208 -1563 2224
rect -1597 1416 -1563 1432
rect -1439 2208 -1405 2224
rect -1439 1416 -1405 1432
rect -1281 2208 -1247 2224
rect -1281 1416 -1247 1432
rect -1123 2208 -1089 2224
rect -1123 1416 -1089 1432
rect -965 2208 -931 2224
rect -965 1416 -931 1432
rect -807 2208 -773 2224
rect -807 1416 -773 1432
rect -649 2208 -615 2224
rect -649 1416 -615 1432
rect -491 2208 -457 2224
rect -491 1416 -457 1432
rect -333 2208 -299 2224
rect -333 1416 -299 1432
rect -175 2208 -141 2224
rect -175 1416 -141 1432
rect -17 2208 17 2224
rect -17 1416 17 1432
rect 141 2208 175 2224
rect 141 1416 175 1432
rect 299 2208 333 2224
rect 299 1416 333 1432
rect 457 2208 491 2224
rect 457 1416 491 1432
rect 615 2208 649 2224
rect 615 1416 649 1432
rect 773 2208 807 2224
rect 773 1416 807 1432
rect 931 2208 965 2224
rect 931 1416 965 1432
rect 1089 2208 1123 2224
rect 1089 1416 1123 1432
rect 1247 2208 1281 2224
rect 1247 1416 1281 1432
rect 1405 2208 1439 2224
rect 1405 1416 1439 1432
rect 1563 2208 1597 2224
rect 1563 1416 1597 1432
rect 1721 2208 1755 2224
rect 1721 1416 1755 1432
rect 1879 2208 1913 2224
rect 1879 1416 1913 1432
rect 2037 2208 2071 2224
rect 2037 1416 2071 1432
rect 2195 2208 2229 2224
rect 2195 1416 2229 1432
rect 2353 2208 2387 2224
rect 2353 1416 2387 1432
rect 2511 2208 2545 2224
rect 2511 1416 2545 1432
rect 2669 2208 2703 2224
rect 2669 1416 2703 1432
rect 2827 2208 2861 2224
rect 2827 1416 2861 1432
rect 2985 2208 3019 2224
rect 2985 1416 3019 1432
rect 3143 2208 3177 2224
rect 3143 1416 3177 1432
rect 3301 2208 3335 2224
rect 3301 1416 3335 1432
rect 3459 2208 3493 2224
rect 3459 1416 3493 1432
rect 3617 2208 3651 2224
rect 3617 1416 3651 1432
rect 3775 2208 3809 2224
rect 3775 1416 3809 1432
rect 3933 2208 3967 2224
rect 3933 1416 3967 1432
rect 4091 2208 4125 2224
rect 4091 1416 4125 1432
rect 4249 2208 4283 2224
rect 4249 1416 4283 1432
rect 4407 2208 4441 2224
rect 4407 1416 4441 1432
rect 4565 2208 4599 2224
rect 4565 1416 4599 1432
rect 4723 2208 4757 2224
rect 4723 1416 4757 1432
rect 4881 2208 4915 2224
rect 4881 1416 4915 1432
rect 5039 2208 5073 2224
rect 5039 1416 5073 1432
rect 5197 2208 5231 2224
rect 5197 1416 5231 1432
rect 5355 2208 5389 2224
rect 5355 1416 5389 1432
rect 5513 2208 5547 2224
rect 5513 1416 5547 1432
rect 5671 2208 5705 2224
rect 5671 1416 5705 1432
rect 5829 2208 5863 2224
rect 5829 1416 5863 1432
rect 5987 2208 6021 2224
rect 5987 1416 6021 1432
rect 6145 2208 6179 2224
rect 6145 1416 6179 1432
rect 6303 2208 6337 2224
rect 6303 1416 6337 1432
rect -6291 1348 -6275 1382
rect -6207 1348 -6191 1382
rect -6133 1348 -6117 1382
rect -6049 1348 -6033 1382
rect -5975 1348 -5959 1382
rect -5891 1348 -5875 1382
rect -5817 1348 -5801 1382
rect -5733 1348 -5717 1382
rect -5659 1348 -5643 1382
rect -5575 1348 -5559 1382
rect -5501 1348 -5485 1382
rect -5417 1348 -5401 1382
rect -5343 1348 -5327 1382
rect -5259 1348 -5243 1382
rect -5185 1348 -5169 1382
rect -5101 1348 -5085 1382
rect -5027 1348 -5011 1382
rect -4943 1348 -4927 1382
rect -4869 1348 -4853 1382
rect -4785 1348 -4769 1382
rect -4711 1348 -4695 1382
rect -4627 1348 -4611 1382
rect -4553 1348 -4537 1382
rect -4469 1348 -4453 1382
rect -4395 1348 -4379 1382
rect -4311 1348 -4295 1382
rect -4237 1348 -4221 1382
rect -4153 1348 -4137 1382
rect -4079 1348 -4063 1382
rect -3995 1348 -3979 1382
rect -3921 1348 -3905 1382
rect -3837 1348 -3821 1382
rect -3763 1348 -3747 1382
rect -3679 1348 -3663 1382
rect -3605 1348 -3589 1382
rect -3521 1348 -3505 1382
rect -3447 1348 -3431 1382
rect -3363 1348 -3347 1382
rect -3289 1348 -3273 1382
rect -3205 1348 -3189 1382
rect -3131 1348 -3115 1382
rect -3047 1348 -3031 1382
rect -2973 1348 -2957 1382
rect -2889 1348 -2873 1382
rect -2815 1348 -2799 1382
rect -2731 1348 -2715 1382
rect -2657 1348 -2641 1382
rect -2573 1348 -2557 1382
rect -2499 1348 -2483 1382
rect -2415 1348 -2399 1382
rect -2341 1348 -2325 1382
rect -2257 1348 -2241 1382
rect -2183 1348 -2167 1382
rect -2099 1348 -2083 1382
rect -2025 1348 -2009 1382
rect -1941 1348 -1925 1382
rect -1867 1348 -1851 1382
rect -1783 1348 -1767 1382
rect -1709 1348 -1693 1382
rect -1625 1348 -1609 1382
rect -1551 1348 -1535 1382
rect -1467 1348 -1451 1382
rect -1393 1348 -1377 1382
rect -1309 1348 -1293 1382
rect -1235 1348 -1219 1382
rect -1151 1348 -1135 1382
rect -1077 1348 -1061 1382
rect -993 1348 -977 1382
rect -919 1348 -903 1382
rect -835 1348 -819 1382
rect -761 1348 -745 1382
rect -677 1348 -661 1382
rect -603 1348 -587 1382
rect -519 1348 -503 1382
rect -445 1348 -429 1382
rect -361 1348 -345 1382
rect -287 1348 -271 1382
rect -203 1348 -187 1382
rect -129 1348 -113 1382
rect -45 1348 -29 1382
rect 29 1348 45 1382
rect 113 1348 129 1382
rect 187 1348 203 1382
rect 271 1348 287 1382
rect 345 1348 361 1382
rect 429 1348 445 1382
rect 503 1348 519 1382
rect 587 1348 603 1382
rect 661 1348 677 1382
rect 745 1348 761 1382
rect 819 1348 835 1382
rect 903 1348 919 1382
rect 977 1348 993 1382
rect 1061 1348 1077 1382
rect 1135 1348 1151 1382
rect 1219 1348 1235 1382
rect 1293 1348 1309 1382
rect 1377 1348 1393 1382
rect 1451 1348 1467 1382
rect 1535 1348 1551 1382
rect 1609 1348 1625 1382
rect 1693 1348 1709 1382
rect 1767 1348 1783 1382
rect 1851 1348 1867 1382
rect 1925 1348 1941 1382
rect 2009 1348 2025 1382
rect 2083 1348 2099 1382
rect 2167 1348 2183 1382
rect 2241 1348 2257 1382
rect 2325 1348 2341 1382
rect 2399 1348 2415 1382
rect 2483 1348 2499 1382
rect 2557 1348 2573 1382
rect 2641 1348 2657 1382
rect 2715 1348 2731 1382
rect 2799 1348 2815 1382
rect 2873 1348 2889 1382
rect 2957 1348 2973 1382
rect 3031 1348 3047 1382
rect 3115 1348 3131 1382
rect 3189 1348 3205 1382
rect 3273 1348 3289 1382
rect 3347 1348 3363 1382
rect 3431 1348 3447 1382
rect 3505 1348 3521 1382
rect 3589 1348 3605 1382
rect 3663 1348 3679 1382
rect 3747 1348 3763 1382
rect 3821 1348 3837 1382
rect 3905 1348 3921 1382
rect 3979 1348 3995 1382
rect 4063 1348 4079 1382
rect 4137 1348 4153 1382
rect 4221 1348 4237 1382
rect 4295 1348 4311 1382
rect 4379 1348 4395 1382
rect 4453 1348 4469 1382
rect 4537 1348 4553 1382
rect 4611 1348 4627 1382
rect 4695 1348 4711 1382
rect 4769 1348 4785 1382
rect 4853 1348 4869 1382
rect 4927 1348 4943 1382
rect 5011 1348 5027 1382
rect 5085 1348 5101 1382
rect 5169 1348 5185 1382
rect 5243 1348 5259 1382
rect 5327 1348 5343 1382
rect 5401 1348 5417 1382
rect 5485 1348 5501 1382
rect 5559 1348 5575 1382
rect 5643 1348 5659 1382
rect 5717 1348 5733 1382
rect 5801 1348 5817 1382
rect 5875 1348 5891 1382
rect 5959 1348 5975 1382
rect 6033 1348 6049 1382
rect 6117 1348 6133 1382
rect 6191 1348 6207 1382
rect 6275 1348 6291 1382
rect -6337 1298 -6303 1314
rect -6337 506 -6303 522
rect -6179 1298 -6145 1314
rect -6179 506 -6145 522
rect -6021 1298 -5987 1314
rect -6021 506 -5987 522
rect -5863 1298 -5829 1314
rect -5863 506 -5829 522
rect -5705 1298 -5671 1314
rect -5705 506 -5671 522
rect -5547 1298 -5513 1314
rect -5547 506 -5513 522
rect -5389 1298 -5355 1314
rect -5389 506 -5355 522
rect -5231 1298 -5197 1314
rect -5231 506 -5197 522
rect -5073 1298 -5039 1314
rect -5073 506 -5039 522
rect -4915 1298 -4881 1314
rect -4915 506 -4881 522
rect -4757 1298 -4723 1314
rect -4757 506 -4723 522
rect -4599 1298 -4565 1314
rect -4599 506 -4565 522
rect -4441 1298 -4407 1314
rect -4441 506 -4407 522
rect -4283 1298 -4249 1314
rect -4283 506 -4249 522
rect -4125 1298 -4091 1314
rect -4125 506 -4091 522
rect -3967 1298 -3933 1314
rect -3967 506 -3933 522
rect -3809 1298 -3775 1314
rect -3809 506 -3775 522
rect -3651 1298 -3617 1314
rect -3651 506 -3617 522
rect -3493 1298 -3459 1314
rect -3493 506 -3459 522
rect -3335 1298 -3301 1314
rect -3335 506 -3301 522
rect -3177 1298 -3143 1314
rect -3177 506 -3143 522
rect -3019 1298 -2985 1314
rect -3019 506 -2985 522
rect -2861 1298 -2827 1314
rect -2861 506 -2827 522
rect -2703 1298 -2669 1314
rect -2703 506 -2669 522
rect -2545 1298 -2511 1314
rect -2545 506 -2511 522
rect -2387 1298 -2353 1314
rect -2387 506 -2353 522
rect -2229 1298 -2195 1314
rect -2229 506 -2195 522
rect -2071 1298 -2037 1314
rect -2071 506 -2037 522
rect -1913 1298 -1879 1314
rect -1913 506 -1879 522
rect -1755 1298 -1721 1314
rect -1755 506 -1721 522
rect -1597 1298 -1563 1314
rect -1597 506 -1563 522
rect -1439 1298 -1405 1314
rect -1439 506 -1405 522
rect -1281 1298 -1247 1314
rect -1281 506 -1247 522
rect -1123 1298 -1089 1314
rect -1123 506 -1089 522
rect -965 1298 -931 1314
rect -965 506 -931 522
rect -807 1298 -773 1314
rect -807 506 -773 522
rect -649 1298 -615 1314
rect -649 506 -615 522
rect -491 1298 -457 1314
rect -491 506 -457 522
rect -333 1298 -299 1314
rect -333 506 -299 522
rect -175 1298 -141 1314
rect -175 506 -141 522
rect -17 1298 17 1314
rect -17 506 17 522
rect 141 1298 175 1314
rect 141 506 175 522
rect 299 1298 333 1314
rect 299 506 333 522
rect 457 1298 491 1314
rect 457 506 491 522
rect 615 1298 649 1314
rect 615 506 649 522
rect 773 1298 807 1314
rect 773 506 807 522
rect 931 1298 965 1314
rect 931 506 965 522
rect 1089 1298 1123 1314
rect 1089 506 1123 522
rect 1247 1298 1281 1314
rect 1247 506 1281 522
rect 1405 1298 1439 1314
rect 1405 506 1439 522
rect 1563 1298 1597 1314
rect 1563 506 1597 522
rect 1721 1298 1755 1314
rect 1721 506 1755 522
rect 1879 1298 1913 1314
rect 1879 506 1913 522
rect 2037 1298 2071 1314
rect 2037 506 2071 522
rect 2195 1298 2229 1314
rect 2195 506 2229 522
rect 2353 1298 2387 1314
rect 2353 506 2387 522
rect 2511 1298 2545 1314
rect 2511 506 2545 522
rect 2669 1298 2703 1314
rect 2669 506 2703 522
rect 2827 1298 2861 1314
rect 2827 506 2861 522
rect 2985 1298 3019 1314
rect 2985 506 3019 522
rect 3143 1298 3177 1314
rect 3143 506 3177 522
rect 3301 1298 3335 1314
rect 3301 506 3335 522
rect 3459 1298 3493 1314
rect 3459 506 3493 522
rect 3617 1298 3651 1314
rect 3617 506 3651 522
rect 3775 1298 3809 1314
rect 3775 506 3809 522
rect 3933 1298 3967 1314
rect 3933 506 3967 522
rect 4091 1298 4125 1314
rect 4091 506 4125 522
rect 4249 1298 4283 1314
rect 4249 506 4283 522
rect 4407 1298 4441 1314
rect 4407 506 4441 522
rect 4565 1298 4599 1314
rect 4565 506 4599 522
rect 4723 1298 4757 1314
rect 4723 506 4757 522
rect 4881 1298 4915 1314
rect 4881 506 4915 522
rect 5039 1298 5073 1314
rect 5039 506 5073 522
rect 5197 1298 5231 1314
rect 5197 506 5231 522
rect 5355 1298 5389 1314
rect 5355 506 5389 522
rect 5513 1298 5547 1314
rect 5513 506 5547 522
rect 5671 1298 5705 1314
rect 5671 506 5705 522
rect 5829 1298 5863 1314
rect 5829 506 5863 522
rect 5987 1298 6021 1314
rect 5987 506 6021 522
rect 6145 1298 6179 1314
rect 6145 506 6179 522
rect 6303 1298 6337 1314
rect 6303 506 6337 522
rect -6291 438 -6275 472
rect -6207 438 -6191 472
rect -6133 438 -6117 472
rect -6049 438 -6033 472
rect -5975 438 -5959 472
rect -5891 438 -5875 472
rect -5817 438 -5801 472
rect -5733 438 -5717 472
rect -5659 438 -5643 472
rect -5575 438 -5559 472
rect -5501 438 -5485 472
rect -5417 438 -5401 472
rect -5343 438 -5327 472
rect -5259 438 -5243 472
rect -5185 438 -5169 472
rect -5101 438 -5085 472
rect -5027 438 -5011 472
rect -4943 438 -4927 472
rect -4869 438 -4853 472
rect -4785 438 -4769 472
rect -4711 438 -4695 472
rect -4627 438 -4611 472
rect -4553 438 -4537 472
rect -4469 438 -4453 472
rect -4395 438 -4379 472
rect -4311 438 -4295 472
rect -4237 438 -4221 472
rect -4153 438 -4137 472
rect -4079 438 -4063 472
rect -3995 438 -3979 472
rect -3921 438 -3905 472
rect -3837 438 -3821 472
rect -3763 438 -3747 472
rect -3679 438 -3663 472
rect -3605 438 -3589 472
rect -3521 438 -3505 472
rect -3447 438 -3431 472
rect -3363 438 -3347 472
rect -3289 438 -3273 472
rect -3205 438 -3189 472
rect -3131 438 -3115 472
rect -3047 438 -3031 472
rect -2973 438 -2957 472
rect -2889 438 -2873 472
rect -2815 438 -2799 472
rect -2731 438 -2715 472
rect -2657 438 -2641 472
rect -2573 438 -2557 472
rect -2499 438 -2483 472
rect -2415 438 -2399 472
rect -2341 438 -2325 472
rect -2257 438 -2241 472
rect -2183 438 -2167 472
rect -2099 438 -2083 472
rect -2025 438 -2009 472
rect -1941 438 -1925 472
rect -1867 438 -1851 472
rect -1783 438 -1767 472
rect -1709 438 -1693 472
rect -1625 438 -1609 472
rect -1551 438 -1535 472
rect -1467 438 -1451 472
rect -1393 438 -1377 472
rect -1309 438 -1293 472
rect -1235 438 -1219 472
rect -1151 438 -1135 472
rect -1077 438 -1061 472
rect -993 438 -977 472
rect -919 438 -903 472
rect -835 438 -819 472
rect -761 438 -745 472
rect -677 438 -661 472
rect -603 438 -587 472
rect -519 438 -503 472
rect -445 438 -429 472
rect -361 438 -345 472
rect -287 438 -271 472
rect -203 438 -187 472
rect -129 438 -113 472
rect -45 438 -29 472
rect 29 438 45 472
rect 113 438 129 472
rect 187 438 203 472
rect 271 438 287 472
rect 345 438 361 472
rect 429 438 445 472
rect 503 438 519 472
rect 587 438 603 472
rect 661 438 677 472
rect 745 438 761 472
rect 819 438 835 472
rect 903 438 919 472
rect 977 438 993 472
rect 1061 438 1077 472
rect 1135 438 1151 472
rect 1219 438 1235 472
rect 1293 438 1309 472
rect 1377 438 1393 472
rect 1451 438 1467 472
rect 1535 438 1551 472
rect 1609 438 1625 472
rect 1693 438 1709 472
rect 1767 438 1783 472
rect 1851 438 1867 472
rect 1925 438 1941 472
rect 2009 438 2025 472
rect 2083 438 2099 472
rect 2167 438 2183 472
rect 2241 438 2257 472
rect 2325 438 2341 472
rect 2399 438 2415 472
rect 2483 438 2499 472
rect 2557 438 2573 472
rect 2641 438 2657 472
rect 2715 438 2731 472
rect 2799 438 2815 472
rect 2873 438 2889 472
rect 2957 438 2973 472
rect 3031 438 3047 472
rect 3115 438 3131 472
rect 3189 438 3205 472
rect 3273 438 3289 472
rect 3347 438 3363 472
rect 3431 438 3447 472
rect 3505 438 3521 472
rect 3589 438 3605 472
rect 3663 438 3679 472
rect 3747 438 3763 472
rect 3821 438 3837 472
rect 3905 438 3921 472
rect 3979 438 3995 472
rect 4063 438 4079 472
rect 4137 438 4153 472
rect 4221 438 4237 472
rect 4295 438 4311 472
rect 4379 438 4395 472
rect 4453 438 4469 472
rect 4537 438 4553 472
rect 4611 438 4627 472
rect 4695 438 4711 472
rect 4769 438 4785 472
rect 4853 438 4869 472
rect 4927 438 4943 472
rect 5011 438 5027 472
rect 5085 438 5101 472
rect 5169 438 5185 472
rect 5243 438 5259 472
rect 5327 438 5343 472
rect 5401 438 5417 472
rect 5485 438 5501 472
rect 5559 438 5575 472
rect 5643 438 5659 472
rect 5717 438 5733 472
rect 5801 438 5817 472
rect 5875 438 5891 472
rect 5959 438 5975 472
rect 6033 438 6049 472
rect 6117 438 6133 472
rect 6191 438 6207 472
rect 6275 438 6291 472
rect -6337 388 -6303 404
rect -6337 -404 -6303 -388
rect -6179 388 -6145 404
rect -6179 -404 -6145 -388
rect -6021 388 -5987 404
rect -6021 -404 -5987 -388
rect -5863 388 -5829 404
rect -5863 -404 -5829 -388
rect -5705 388 -5671 404
rect -5705 -404 -5671 -388
rect -5547 388 -5513 404
rect -5547 -404 -5513 -388
rect -5389 388 -5355 404
rect -5389 -404 -5355 -388
rect -5231 388 -5197 404
rect -5231 -404 -5197 -388
rect -5073 388 -5039 404
rect -5073 -404 -5039 -388
rect -4915 388 -4881 404
rect -4915 -404 -4881 -388
rect -4757 388 -4723 404
rect -4757 -404 -4723 -388
rect -4599 388 -4565 404
rect -4599 -404 -4565 -388
rect -4441 388 -4407 404
rect -4441 -404 -4407 -388
rect -4283 388 -4249 404
rect -4283 -404 -4249 -388
rect -4125 388 -4091 404
rect -4125 -404 -4091 -388
rect -3967 388 -3933 404
rect -3967 -404 -3933 -388
rect -3809 388 -3775 404
rect -3809 -404 -3775 -388
rect -3651 388 -3617 404
rect -3651 -404 -3617 -388
rect -3493 388 -3459 404
rect -3493 -404 -3459 -388
rect -3335 388 -3301 404
rect -3335 -404 -3301 -388
rect -3177 388 -3143 404
rect -3177 -404 -3143 -388
rect -3019 388 -2985 404
rect -3019 -404 -2985 -388
rect -2861 388 -2827 404
rect -2861 -404 -2827 -388
rect -2703 388 -2669 404
rect -2703 -404 -2669 -388
rect -2545 388 -2511 404
rect -2545 -404 -2511 -388
rect -2387 388 -2353 404
rect -2387 -404 -2353 -388
rect -2229 388 -2195 404
rect -2229 -404 -2195 -388
rect -2071 388 -2037 404
rect -2071 -404 -2037 -388
rect -1913 388 -1879 404
rect -1913 -404 -1879 -388
rect -1755 388 -1721 404
rect -1755 -404 -1721 -388
rect -1597 388 -1563 404
rect -1597 -404 -1563 -388
rect -1439 388 -1405 404
rect -1439 -404 -1405 -388
rect -1281 388 -1247 404
rect -1281 -404 -1247 -388
rect -1123 388 -1089 404
rect -1123 -404 -1089 -388
rect -965 388 -931 404
rect -965 -404 -931 -388
rect -807 388 -773 404
rect -807 -404 -773 -388
rect -649 388 -615 404
rect -649 -404 -615 -388
rect -491 388 -457 404
rect -491 -404 -457 -388
rect -333 388 -299 404
rect -333 -404 -299 -388
rect -175 388 -141 404
rect -175 -404 -141 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 141 388 175 404
rect 141 -404 175 -388
rect 299 388 333 404
rect 299 -404 333 -388
rect 457 388 491 404
rect 457 -404 491 -388
rect 615 388 649 404
rect 615 -404 649 -388
rect 773 388 807 404
rect 773 -404 807 -388
rect 931 388 965 404
rect 931 -404 965 -388
rect 1089 388 1123 404
rect 1089 -404 1123 -388
rect 1247 388 1281 404
rect 1247 -404 1281 -388
rect 1405 388 1439 404
rect 1405 -404 1439 -388
rect 1563 388 1597 404
rect 1563 -404 1597 -388
rect 1721 388 1755 404
rect 1721 -404 1755 -388
rect 1879 388 1913 404
rect 1879 -404 1913 -388
rect 2037 388 2071 404
rect 2037 -404 2071 -388
rect 2195 388 2229 404
rect 2195 -404 2229 -388
rect 2353 388 2387 404
rect 2353 -404 2387 -388
rect 2511 388 2545 404
rect 2511 -404 2545 -388
rect 2669 388 2703 404
rect 2669 -404 2703 -388
rect 2827 388 2861 404
rect 2827 -404 2861 -388
rect 2985 388 3019 404
rect 2985 -404 3019 -388
rect 3143 388 3177 404
rect 3143 -404 3177 -388
rect 3301 388 3335 404
rect 3301 -404 3335 -388
rect 3459 388 3493 404
rect 3459 -404 3493 -388
rect 3617 388 3651 404
rect 3617 -404 3651 -388
rect 3775 388 3809 404
rect 3775 -404 3809 -388
rect 3933 388 3967 404
rect 3933 -404 3967 -388
rect 4091 388 4125 404
rect 4091 -404 4125 -388
rect 4249 388 4283 404
rect 4249 -404 4283 -388
rect 4407 388 4441 404
rect 4407 -404 4441 -388
rect 4565 388 4599 404
rect 4565 -404 4599 -388
rect 4723 388 4757 404
rect 4723 -404 4757 -388
rect 4881 388 4915 404
rect 4881 -404 4915 -388
rect 5039 388 5073 404
rect 5039 -404 5073 -388
rect 5197 388 5231 404
rect 5197 -404 5231 -388
rect 5355 388 5389 404
rect 5355 -404 5389 -388
rect 5513 388 5547 404
rect 5513 -404 5547 -388
rect 5671 388 5705 404
rect 5671 -404 5705 -388
rect 5829 388 5863 404
rect 5829 -404 5863 -388
rect 5987 388 6021 404
rect 5987 -404 6021 -388
rect 6145 388 6179 404
rect 6145 -404 6179 -388
rect 6303 388 6337 404
rect 6303 -404 6337 -388
rect -6291 -472 -6275 -438
rect -6207 -472 -6191 -438
rect -6133 -472 -6117 -438
rect -6049 -472 -6033 -438
rect -5975 -472 -5959 -438
rect -5891 -472 -5875 -438
rect -5817 -472 -5801 -438
rect -5733 -472 -5717 -438
rect -5659 -472 -5643 -438
rect -5575 -472 -5559 -438
rect -5501 -472 -5485 -438
rect -5417 -472 -5401 -438
rect -5343 -472 -5327 -438
rect -5259 -472 -5243 -438
rect -5185 -472 -5169 -438
rect -5101 -472 -5085 -438
rect -5027 -472 -5011 -438
rect -4943 -472 -4927 -438
rect -4869 -472 -4853 -438
rect -4785 -472 -4769 -438
rect -4711 -472 -4695 -438
rect -4627 -472 -4611 -438
rect -4553 -472 -4537 -438
rect -4469 -472 -4453 -438
rect -4395 -472 -4379 -438
rect -4311 -472 -4295 -438
rect -4237 -472 -4221 -438
rect -4153 -472 -4137 -438
rect -4079 -472 -4063 -438
rect -3995 -472 -3979 -438
rect -3921 -472 -3905 -438
rect -3837 -472 -3821 -438
rect -3763 -472 -3747 -438
rect -3679 -472 -3663 -438
rect -3605 -472 -3589 -438
rect -3521 -472 -3505 -438
rect -3447 -472 -3431 -438
rect -3363 -472 -3347 -438
rect -3289 -472 -3273 -438
rect -3205 -472 -3189 -438
rect -3131 -472 -3115 -438
rect -3047 -472 -3031 -438
rect -2973 -472 -2957 -438
rect -2889 -472 -2873 -438
rect -2815 -472 -2799 -438
rect -2731 -472 -2715 -438
rect -2657 -472 -2641 -438
rect -2573 -472 -2557 -438
rect -2499 -472 -2483 -438
rect -2415 -472 -2399 -438
rect -2341 -472 -2325 -438
rect -2257 -472 -2241 -438
rect -2183 -472 -2167 -438
rect -2099 -472 -2083 -438
rect -2025 -472 -2009 -438
rect -1941 -472 -1925 -438
rect -1867 -472 -1851 -438
rect -1783 -472 -1767 -438
rect -1709 -472 -1693 -438
rect -1625 -472 -1609 -438
rect -1551 -472 -1535 -438
rect -1467 -472 -1451 -438
rect -1393 -472 -1377 -438
rect -1309 -472 -1293 -438
rect -1235 -472 -1219 -438
rect -1151 -472 -1135 -438
rect -1077 -472 -1061 -438
rect -993 -472 -977 -438
rect -919 -472 -903 -438
rect -835 -472 -819 -438
rect -761 -472 -745 -438
rect -677 -472 -661 -438
rect -603 -472 -587 -438
rect -519 -472 -503 -438
rect -445 -472 -429 -438
rect -361 -472 -345 -438
rect -287 -472 -271 -438
rect -203 -472 -187 -438
rect -129 -472 -113 -438
rect -45 -472 -29 -438
rect 29 -472 45 -438
rect 113 -472 129 -438
rect 187 -472 203 -438
rect 271 -472 287 -438
rect 345 -472 361 -438
rect 429 -472 445 -438
rect 503 -472 519 -438
rect 587 -472 603 -438
rect 661 -472 677 -438
rect 745 -472 761 -438
rect 819 -472 835 -438
rect 903 -472 919 -438
rect 977 -472 993 -438
rect 1061 -472 1077 -438
rect 1135 -472 1151 -438
rect 1219 -472 1235 -438
rect 1293 -472 1309 -438
rect 1377 -472 1393 -438
rect 1451 -472 1467 -438
rect 1535 -472 1551 -438
rect 1609 -472 1625 -438
rect 1693 -472 1709 -438
rect 1767 -472 1783 -438
rect 1851 -472 1867 -438
rect 1925 -472 1941 -438
rect 2009 -472 2025 -438
rect 2083 -472 2099 -438
rect 2167 -472 2183 -438
rect 2241 -472 2257 -438
rect 2325 -472 2341 -438
rect 2399 -472 2415 -438
rect 2483 -472 2499 -438
rect 2557 -472 2573 -438
rect 2641 -472 2657 -438
rect 2715 -472 2731 -438
rect 2799 -472 2815 -438
rect 2873 -472 2889 -438
rect 2957 -472 2973 -438
rect 3031 -472 3047 -438
rect 3115 -472 3131 -438
rect 3189 -472 3205 -438
rect 3273 -472 3289 -438
rect 3347 -472 3363 -438
rect 3431 -472 3447 -438
rect 3505 -472 3521 -438
rect 3589 -472 3605 -438
rect 3663 -472 3679 -438
rect 3747 -472 3763 -438
rect 3821 -472 3837 -438
rect 3905 -472 3921 -438
rect 3979 -472 3995 -438
rect 4063 -472 4079 -438
rect 4137 -472 4153 -438
rect 4221 -472 4237 -438
rect 4295 -472 4311 -438
rect 4379 -472 4395 -438
rect 4453 -472 4469 -438
rect 4537 -472 4553 -438
rect 4611 -472 4627 -438
rect 4695 -472 4711 -438
rect 4769 -472 4785 -438
rect 4853 -472 4869 -438
rect 4927 -472 4943 -438
rect 5011 -472 5027 -438
rect 5085 -472 5101 -438
rect 5169 -472 5185 -438
rect 5243 -472 5259 -438
rect 5327 -472 5343 -438
rect 5401 -472 5417 -438
rect 5485 -472 5501 -438
rect 5559 -472 5575 -438
rect 5643 -472 5659 -438
rect 5717 -472 5733 -438
rect 5801 -472 5817 -438
rect 5875 -472 5891 -438
rect 5959 -472 5975 -438
rect 6033 -472 6049 -438
rect 6117 -472 6133 -438
rect 6191 -472 6207 -438
rect 6275 -472 6291 -438
rect -6337 -522 -6303 -506
rect -6337 -1314 -6303 -1298
rect -6179 -522 -6145 -506
rect -6179 -1314 -6145 -1298
rect -6021 -522 -5987 -506
rect -6021 -1314 -5987 -1298
rect -5863 -522 -5829 -506
rect -5863 -1314 -5829 -1298
rect -5705 -522 -5671 -506
rect -5705 -1314 -5671 -1298
rect -5547 -522 -5513 -506
rect -5547 -1314 -5513 -1298
rect -5389 -522 -5355 -506
rect -5389 -1314 -5355 -1298
rect -5231 -522 -5197 -506
rect -5231 -1314 -5197 -1298
rect -5073 -522 -5039 -506
rect -5073 -1314 -5039 -1298
rect -4915 -522 -4881 -506
rect -4915 -1314 -4881 -1298
rect -4757 -522 -4723 -506
rect -4757 -1314 -4723 -1298
rect -4599 -522 -4565 -506
rect -4599 -1314 -4565 -1298
rect -4441 -522 -4407 -506
rect -4441 -1314 -4407 -1298
rect -4283 -522 -4249 -506
rect -4283 -1314 -4249 -1298
rect -4125 -522 -4091 -506
rect -4125 -1314 -4091 -1298
rect -3967 -522 -3933 -506
rect -3967 -1314 -3933 -1298
rect -3809 -522 -3775 -506
rect -3809 -1314 -3775 -1298
rect -3651 -522 -3617 -506
rect -3651 -1314 -3617 -1298
rect -3493 -522 -3459 -506
rect -3493 -1314 -3459 -1298
rect -3335 -522 -3301 -506
rect -3335 -1314 -3301 -1298
rect -3177 -522 -3143 -506
rect -3177 -1314 -3143 -1298
rect -3019 -522 -2985 -506
rect -3019 -1314 -2985 -1298
rect -2861 -522 -2827 -506
rect -2861 -1314 -2827 -1298
rect -2703 -522 -2669 -506
rect -2703 -1314 -2669 -1298
rect -2545 -522 -2511 -506
rect -2545 -1314 -2511 -1298
rect -2387 -522 -2353 -506
rect -2387 -1314 -2353 -1298
rect -2229 -522 -2195 -506
rect -2229 -1314 -2195 -1298
rect -2071 -522 -2037 -506
rect -2071 -1314 -2037 -1298
rect -1913 -522 -1879 -506
rect -1913 -1314 -1879 -1298
rect -1755 -522 -1721 -506
rect -1755 -1314 -1721 -1298
rect -1597 -522 -1563 -506
rect -1597 -1314 -1563 -1298
rect -1439 -522 -1405 -506
rect -1439 -1314 -1405 -1298
rect -1281 -522 -1247 -506
rect -1281 -1314 -1247 -1298
rect -1123 -522 -1089 -506
rect -1123 -1314 -1089 -1298
rect -965 -522 -931 -506
rect -965 -1314 -931 -1298
rect -807 -522 -773 -506
rect -807 -1314 -773 -1298
rect -649 -522 -615 -506
rect -649 -1314 -615 -1298
rect -491 -522 -457 -506
rect -491 -1314 -457 -1298
rect -333 -522 -299 -506
rect -333 -1314 -299 -1298
rect -175 -522 -141 -506
rect -175 -1314 -141 -1298
rect -17 -522 17 -506
rect -17 -1314 17 -1298
rect 141 -522 175 -506
rect 141 -1314 175 -1298
rect 299 -522 333 -506
rect 299 -1314 333 -1298
rect 457 -522 491 -506
rect 457 -1314 491 -1298
rect 615 -522 649 -506
rect 615 -1314 649 -1298
rect 773 -522 807 -506
rect 773 -1314 807 -1298
rect 931 -522 965 -506
rect 931 -1314 965 -1298
rect 1089 -522 1123 -506
rect 1089 -1314 1123 -1298
rect 1247 -522 1281 -506
rect 1247 -1314 1281 -1298
rect 1405 -522 1439 -506
rect 1405 -1314 1439 -1298
rect 1563 -522 1597 -506
rect 1563 -1314 1597 -1298
rect 1721 -522 1755 -506
rect 1721 -1314 1755 -1298
rect 1879 -522 1913 -506
rect 1879 -1314 1913 -1298
rect 2037 -522 2071 -506
rect 2037 -1314 2071 -1298
rect 2195 -522 2229 -506
rect 2195 -1314 2229 -1298
rect 2353 -522 2387 -506
rect 2353 -1314 2387 -1298
rect 2511 -522 2545 -506
rect 2511 -1314 2545 -1298
rect 2669 -522 2703 -506
rect 2669 -1314 2703 -1298
rect 2827 -522 2861 -506
rect 2827 -1314 2861 -1298
rect 2985 -522 3019 -506
rect 2985 -1314 3019 -1298
rect 3143 -522 3177 -506
rect 3143 -1314 3177 -1298
rect 3301 -522 3335 -506
rect 3301 -1314 3335 -1298
rect 3459 -522 3493 -506
rect 3459 -1314 3493 -1298
rect 3617 -522 3651 -506
rect 3617 -1314 3651 -1298
rect 3775 -522 3809 -506
rect 3775 -1314 3809 -1298
rect 3933 -522 3967 -506
rect 3933 -1314 3967 -1298
rect 4091 -522 4125 -506
rect 4091 -1314 4125 -1298
rect 4249 -522 4283 -506
rect 4249 -1314 4283 -1298
rect 4407 -522 4441 -506
rect 4407 -1314 4441 -1298
rect 4565 -522 4599 -506
rect 4565 -1314 4599 -1298
rect 4723 -522 4757 -506
rect 4723 -1314 4757 -1298
rect 4881 -522 4915 -506
rect 4881 -1314 4915 -1298
rect 5039 -522 5073 -506
rect 5039 -1314 5073 -1298
rect 5197 -522 5231 -506
rect 5197 -1314 5231 -1298
rect 5355 -522 5389 -506
rect 5355 -1314 5389 -1298
rect 5513 -522 5547 -506
rect 5513 -1314 5547 -1298
rect 5671 -522 5705 -506
rect 5671 -1314 5705 -1298
rect 5829 -522 5863 -506
rect 5829 -1314 5863 -1298
rect 5987 -522 6021 -506
rect 5987 -1314 6021 -1298
rect 6145 -522 6179 -506
rect 6145 -1314 6179 -1298
rect 6303 -522 6337 -506
rect 6303 -1314 6337 -1298
rect -6291 -1382 -6275 -1348
rect -6207 -1382 -6191 -1348
rect -6133 -1382 -6117 -1348
rect -6049 -1382 -6033 -1348
rect -5975 -1382 -5959 -1348
rect -5891 -1382 -5875 -1348
rect -5817 -1382 -5801 -1348
rect -5733 -1382 -5717 -1348
rect -5659 -1382 -5643 -1348
rect -5575 -1382 -5559 -1348
rect -5501 -1382 -5485 -1348
rect -5417 -1382 -5401 -1348
rect -5343 -1382 -5327 -1348
rect -5259 -1382 -5243 -1348
rect -5185 -1382 -5169 -1348
rect -5101 -1382 -5085 -1348
rect -5027 -1382 -5011 -1348
rect -4943 -1382 -4927 -1348
rect -4869 -1382 -4853 -1348
rect -4785 -1382 -4769 -1348
rect -4711 -1382 -4695 -1348
rect -4627 -1382 -4611 -1348
rect -4553 -1382 -4537 -1348
rect -4469 -1382 -4453 -1348
rect -4395 -1382 -4379 -1348
rect -4311 -1382 -4295 -1348
rect -4237 -1382 -4221 -1348
rect -4153 -1382 -4137 -1348
rect -4079 -1382 -4063 -1348
rect -3995 -1382 -3979 -1348
rect -3921 -1382 -3905 -1348
rect -3837 -1382 -3821 -1348
rect -3763 -1382 -3747 -1348
rect -3679 -1382 -3663 -1348
rect -3605 -1382 -3589 -1348
rect -3521 -1382 -3505 -1348
rect -3447 -1382 -3431 -1348
rect -3363 -1382 -3347 -1348
rect -3289 -1382 -3273 -1348
rect -3205 -1382 -3189 -1348
rect -3131 -1382 -3115 -1348
rect -3047 -1382 -3031 -1348
rect -2973 -1382 -2957 -1348
rect -2889 -1382 -2873 -1348
rect -2815 -1382 -2799 -1348
rect -2731 -1382 -2715 -1348
rect -2657 -1382 -2641 -1348
rect -2573 -1382 -2557 -1348
rect -2499 -1382 -2483 -1348
rect -2415 -1382 -2399 -1348
rect -2341 -1382 -2325 -1348
rect -2257 -1382 -2241 -1348
rect -2183 -1382 -2167 -1348
rect -2099 -1382 -2083 -1348
rect -2025 -1382 -2009 -1348
rect -1941 -1382 -1925 -1348
rect -1867 -1382 -1851 -1348
rect -1783 -1382 -1767 -1348
rect -1709 -1382 -1693 -1348
rect -1625 -1382 -1609 -1348
rect -1551 -1382 -1535 -1348
rect -1467 -1382 -1451 -1348
rect -1393 -1382 -1377 -1348
rect -1309 -1382 -1293 -1348
rect -1235 -1382 -1219 -1348
rect -1151 -1382 -1135 -1348
rect -1077 -1382 -1061 -1348
rect -993 -1382 -977 -1348
rect -919 -1382 -903 -1348
rect -835 -1382 -819 -1348
rect -761 -1382 -745 -1348
rect -677 -1382 -661 -1348
rect -603 -1382 -587 -1348
rect -519 -1382 -503 -1348
rect -445 -1382 -429 -1348
rect -361 -1382 -345 -1348
rect -287 -1382 -271 -1348
rect -203 -1382 -187 -1348
rect -129 -1382 -113 -1348
rect -45 -1382 -29 -1348
rect 29 -1382 45 -1348
rect 113 -1382 129 -1348
rect 187 -1382 203 -1348
rect 271 -1382 287 -1348
rect 345 -1382 361 -1348
rect 429 -1382 445 -1348
rect 503 -1382 519 -1348
rect 587 -1382 603 -1348
rect 661 -1382 677 -1348
rect 745 -1382 761 -1348
rect 819 -1382 835 -1348
rect 903 -1382 919 -1348
rect 977 -1382 993 -1348
rect 1061 -1382 1077 -1348
rect 1135 -1382 1151 -1348
rect 1219 -1382 1235 -1348
rect 1293 -1382 1309 -1348
rect 1377 -1382 1393 -1348
rect 1451 -1382 1467 -1348
rect 1535 -1382 1551 -1348
rect 1609 -1382 1625 -1348
rect 1693 -1382 1709 -1348
rect 1767 -1382 1783 -1348
rect 1851 -1382 1867 -1348
rect 1925 -1382 1941 -1348
rect 2009 -1382 2025 -1348
rect 2083 -1382 2099 -1348
rect 2167 -1382 2183 -1348
rect 2241 -1382 2257 -1348
rect 2325 -1382 2341 -1348
rect 2399 -1382 2415 -1348
rect 2483 -1382 2499 -1348
rect 2557 -1382 2573 -1348
rect 2641 -1382 2657 -1348
rect 2715 -1382 2731 -1348
rect 2799 -1382 2815 -1348
rect 2873 -1382 2889 -1348
rect 2957 -1382 2973 -1348
rect 3031 -1382 3047 -1348
rect 3115 -1382 3131 -1348
rect 3189 -1382 3205 -1348
rect 3273 -1382 3289 -1348
rect 3347 -1382 3363 -1348
rect 3431 -1382 3447 -1348
rect 3505 -1382 3521 -1348
rect 3589 -1382 3605 -1348
rect 3663 -1382 3679 -1348
rect 3747 -1382 3763 -1348
rect 3821 -1382 3837 -1348
rect 3905 -1382 3921 -1348
rect 3979 -1382 3995 -1348
rect 4063 -1382 4079 -1348
rect 4137 -1382 4153 -1348
rect 4221 -1382 4237 -1348
rect 4295 -1382 4311 -1348
rect 4379 -1382 4395 -1348
rect 4453 -1382 4469 -1348
rect 4537 -1382 4553 -1348
rect 4611 -1382 4627 -1348
rect 4695 -1382 4711 -1348
rect 4769 -1382 4785 -1348
rect 4853 -1382 4869 -1348
rect 4927 -1382 4943 -1348
rect 5011 -1382 5027 -1348
rect 5085 -1382 5101 -1348
rect 5169 -1382 5185 -1348
rect 5243 -1382 5259 -1348
rect 5327 -1382 5343 -1348
rect 5401 -1382 5417 -1348
rect 5485 -1382 5501 -1348
rect 5559 -1382 5575 -1348
rect 5643 -1382 5659 -1348
rect 5717 -1382 5733 -1348
rect 5801 -1382 5817 -1348
rect 5875 -1382 5891 -1348
rect 5959 -1382 5975 -1348
rect 6033 -1382 6049 -1348
rect 6117 -1382 6133 -1348
rect 6191 -1382 6207 -1348
rect 6275 -1382 6291 -1348
rect -6337 -1432 -6303 -1416
rect -6337 -2224 -6303 -2208
rect -6179 -1432 -6145 -1416
rect -6179 -2224 -6145 -2208
rect -6021 -1432 -5987 -1416
rect -6021 -2224 -5987 -2208
rect -5863 -1432 -5829 -1416
rect -5863 -2224 -5829 -2208
rect -5705 -1432 -5671 -1416
rect -5705 -2224 -5671 -2208
rect -5547 -1432 -5513 -1416
rect -5547 -2224 -5513 -2208
rect -5389 -1432 -5355 -1416
rect -5389 -2224 -5355 -2208
rect -5231 -1432 -5197 -1416
rect -5231 -2224 -5197 -2208
rect -5073 -1432 -5039 -1416
rect -5073 -2224 -5039 -2208
rect -4915 -1432 -4881 -1416
rect -4915 -2224 -4881 -2208
rect -4757 -1432 -4723 -1416
rect -4757 -2224 -4723 -2208
rect -4599 -1432 -4565 -1416
rect -4599 -2224 -4565 -2208
rect -4441 -1432 -4407 -1416
rect -4441 -2224 -4407 -2208
rect -4283 -1432 -4249 -1416
rect -4283 -2224 -4249 -2208
rect -4125 -1432 -4091 -1416
rect -4125 -2224 -4091 -2208
rect -3967 -1432 -3933 -1416
rect -3967 -2224 -3933 -2208
rect -3809 -1432 -3775 -1416
rect -3809 -2224 -3775 -2208
rect -3651 -1432 -3617 -1416
rect -3651 -2224 -3617 -2208
rect -3493 -1432 -3459 -1416
rect -3493 -2224 -3459 -2208
rect -3335 -1432 -3301 -1416
rect -3335 -2224 -3301 -2208
rect -3177 -1432 -3143 -1416
rect -3177 -2224 -3143 -2208
rect -3019 -1432 -2985 -1416
rect -3019 -2224 -2985 -2208
rect -2861 -1432 -2827 -1416
rect -2861 -2224 -2827 -2208
rect -2703 -1432 -2669 -1416
rect -2703 -2224 -2669 -2208
rect -2545 -1432 -2511 -1416
rect -2545 -2224 -2511 -2208
rect -2387 -1432 -2353 -1416
rect -2387 -2224 -2353 -2208
rect -2229 -1432 -2195 -1416
rect -2229 -2224 -2195 -2208
rect -2071 -1432 -2037 -1416
rect -2071 -2224 -2037 -2208
rect -1913 -1432 -1879 -1416
rect -1913 -2224 -1879 -2208
rect -1755 -1432 -1721 -1416
rect -1755 -2224 -1721 -2208
rect -1597 -1432 -1563 -1416
rect -1597 -2224 -1563 -2208
rect -1439 -1432 -1405 -1416
rect -1439 -2224 -1405 -2208
rect -1281 -1432 -1247 -1416
rect -1281 -2224 -1247 -2208
rect -1123 -1432 -1089 -1416
rect -1123 -2224 -1089 -2208
rect -965 -1432 -931 -1416
rect -965 -2224 -931 -2208
rect -807 -1432 -773 -1416
rect -807 -2224 -773 -2208
rect -649 -1432 -615 -1416
rect -649 -2224 -615 -2208
rect -491 -1432 -457 -1416
rect -491 -2224 -457 -2208
rect -333 -1432 -299 -1416
rect -333 -2224 -299 -2208
rect -175 -1432 -141 -1416
rect -175 -2224 -141 -2208
rect -17 -1432 17 -1416
rect -17 -2224 17 -2208
rect 141 -1432 175 -1416
rect 141 -2224 175 -2208
rect 299 -1432 333 -1416
rect 299 -2224 333 -2208
rect 457 -1432 491 -1416
rect 457 -2224 491 -2208
rect 615 -1432 649 -1416
rect 615 -2224 649 -2208
rect 773 -1432 807 -1416
rect 773 -2224 807 -2208
rect 931 -1432 965 -1416
rect 931 -2224 965 -2208
rect 1089 -1432 1123 -1416
rect 1089 -2224 1123 -2208
rect 1247 -1432 1281 -1416
rect 1247 -2224 1281 -2208
rect 1405 -1432 1439 -1416
rect 1405 -2224 1439 -2208
rect 1563 -1432 1597 -1416
rect 1563 -2224 1597 -2208
rect 1721 -1432 1755 -1416
rect 1721 -2224 1755 -2208
rect 1879 -1432 1913 -1416
rect 1879 -2224 1913 -2208
rect 2037 -1432 2071 -1416
rect 2037 -2224 2071 -2208
rect 2195 -1432 2229 -1416
rect 2195 -2224 2229 -2208
rect 2353 -1432 2387 -1416
rect 2353 -2224 2387 -2208
rect 2511 -1432 2545 -1416
rect 2511 -2224 2545 -2208
rect 2669 -1432 2703 -1416
rect 2669 -2224 2703 -2208
rect 2827 -1432 2861 -1416
rect 2827 -2224 2861 -2208
rect 2985 -1432 3019 -1416
rect 2985 -2224 3019 -2208
rect 3143 -1432 3177 -1416
rect 3143 -2224 3177 -2208
rect 3301 -1432 3335 -1416
rect 3301 -2224 3335 -2208
rect 3459 -1432 3493 -1416
rect 3459 -2224 3493 -2208
rect 3617 -1432 3651 -1416
rect 3617 -2224 3651 -2208
rect 3775 -1432 3809 -1416
rect 3775 -2224 3809 -2208
rect 3933 -1432 3967 -1416
rect 3933 -2224 3967 -2208
rect 4091 -1432 4125 -1416
rect 4091 -2224 4125 -2208
rect 4249 -1432 4283 -1416
rect 4249 -2224 4283 -2208
rect 4407 -1432 4441 -1416
rect 4407 -2224 4441 -2208
rect 4565 -1432 4599 -1416
rect 4565 -2224 4599 -2208
rect 4723 -1432 4757 -1416
rect 4723 -2224 4757 -2208
rect 4881 -1432 4915 -1416
rect 4881 -2224 4915 -2208
rect 5039 -1432 5073 -1416
rect 5039 -2224 5073 -2208
rect 5197 -1432 5231 -1416
rect 5197 -2224 5231 -2208
rect 5355 -1432 5389 -1416
rect 5355 -2224 5389 -2208
rect 5513 -1432 5547 -1416
rect 5513 -2224 5547 -2208
rect 5671 -1432 5705 -1416
rect 5671 -2224 5705 -2208
rect 5829 -1432 5863 -1416
rect 5829 -2224 5863 -2208
rect 5987 -1432 6021 -1416
rect 5987 -2224 6021 -2208
rect 6145 -1432 6179 -1416
rect 6145 -2224 6179 -2208
rect 6303 -1432 6337 -1416
rect 6303 -2224 6337 -2208
rect -6291 -2292 -6275 -2258
rect -6207 -2292 -6191 -2258
rect -6133 -2292 -6117 -2258
rect -6049 -2292 -6033 -2258
rect -5975 -2292 -5959 -2258
rect -5891 -2292 -5875 -2258
rect -5817 -2292 -5801 -2258
rect -5733 -2292 -5717 -2258
rect -5659 -2292 -5643 -2258
rect -5575 -2292 -5559 -2258
rect -5501 -2292 -5485 -2258
rect -5417 -2292 -5401 -2258
rect -5343 -2292 -5327 -2258
rect -5259 -2292 -5243 -2258
rect -5185 -2292 -5169 -2258
rect -5101 -2292 -5085 -2258
rect -5027 -2292 -5011 -2258
rect -4943 -2292 -4927 -2258
rect -4869 -2292 -4853 -2258
rect -4785 -2292 -4769 -2258
rect -4711 -2292 -4695 -2258
rect -4627 -2292 -4611 -2258
rect -4553 -2292 -4537 -2258
rect -4469 -2292 -4453 -2258
rect -4395 -2292 -4379 -2258
rect -4311 -2292 -4295 -2258
rect -4237 -2292 -4221 -2258
rect -4153 -2292 -4137 -2258
rect -4079 -2292 -4063 -2258
rect -3995 -2292 -3979 -2258
rect -3921 -2292 -3905 -2258
rect -3837 -2292 -3821 -2258
rect -3763 -2292 -3747 -2258
rect -3679 -2292 -3663 -2258
rect -3605 -2292 -3589 -2258
rect -3521 -2292 -3505 -2258
rect -3447 -2292 -3431 -2258
rect -3363 -2292 -3347 -2258
rect -3289 -2292 -3273 -2258
rect -3205 -2292 -3189 -2258
rect -3131 -2292 -3115 -2258
rect -3047 -2292 -3031 -2258
rect -2973 -2292 -2957 -2258
rect -2889 -2292 -2873 -2258
rect -2815 -2292 -2799 -2258
rect -2731 -2292 -2715 -2258
rect -2657 -2292 -2641 -2258
rect -2573 -2292 -2557 -2258
rect -2499 -2292 -2483 -2258
rect -2415 -2292 -2399 -2258
rect -2341 -2292 -2325 -2258
rect -2257 -2292 -2241 -2258
rect -2183 -2292 -2167 -2258
rect -2099 -2292 -2083 -2258
rect -2025 -2292 -2009 -2258
rect -1941 -2292 -1925 -2258
rect -1867 -2292 -1851 -2258
rect -1783 -2292 -1767 -2258
rect -1709 -2292 -1693 -2258
rect -1625 -2292 -1609 -2258
rect -1551 -2292 -1535 -2258
rect -1467 -2292 -1451 -2258
rect -1393 -2292 -1377 -2258
rect -1309 -2292 -1293 -2258
rect -1235 -2292 -1219 -2258
rect -1151 -2292 -1135 -2258
rect -1077 -2292 -1061 -2258
rect -993 -2292 -977 -2258
rect -919 -2292 -903 -2258
rect -835 -2292 -819 -2258
rect -761 -2292 -745 -2258
rect -677 -2292 -661 -2258
rect -603 -2292 -587 -2258
rect -519 -2292 -503 -2258
rect -445 -2292 -429 -2258
rect -361 -2292 -345 -2258
rect -287 -2292 -271 -2258
rect -203 -2292 -187 -2258
rect -129 -2292 -113 -2258
rect -45 -2292 -29 -2258
rect 29 -2292 45 -2258
rect 113 -2292 129 -2258
rect 187 -2292 203 -2258
rect 271 -2292 287 -2258
rect 345 -2292 361 -2258
rect 429 -2292 445 -2258
rect 503 -2292 519 -2258
rect 587 -2292 603 -2258
rect 661 -2292 677 -2258
rect 745 -2292 761 -2258
rect 819 -2292 835 -2258
rect 903 -2292 919 -2258
rect 977 -2292 993 -2258
rect 1061 -2292 1077 -2258
rect 1135 -2292 1151 -2258
rect 1219 -2292 1235 -2258
rect 1293 -2292 1309 -2258
rect 1377 -2292 1393 -2258
rect 1451 -2292 1467 -2258
rect 1535 -2292 1551 -2258
rect 1609 -2292 1625 -2258
rect 1693 -2292 1709 -2258
rect 1767 -2292 1783 -2258
rect 1851 -2292 1867 -2258
rect 1925 -2292 1941 -2258
rect 2009 -2292 2025 -2258
rect 2083 -2292 2099 -2258
rect 2167 -2292 2183 -2258
rect 2241 -2292 2257 -2258
rect 2325 -2292 2341 -2258
rect 2399 -2292 2415 -2258
rect 2483 -2292 2499 -2258
rect 2557 -2292 2573 -2258
rect 2641 -2292 2657 -2258
rect 2715 -2292 2731 -2258
rect 2799 -2292 2815 -2258
rect 2873 -2292 2889 -2258
rect 2957 -2292 2973 -2258
rect 3031 -2292 3047 -2258
rect 3115 -2292 3131 -2258
rect 3189 -2292 3205 -2258
rect 3273 -2292 3289 -2258
rect 3347 -2292 3363 -2258
rect 3431 -2292 3447 -2258
rect 3505 -2292 3521 -2258
rect 3589 -2292 3605 -2258
rect 3663 -2292 3679 -2258
rect 3747 -2292 3763 -2258
rect 3821 -2292 3837 -2258
rect 3905 -2292 3921 -2258
rect 3979 -2292 3995 -2258
rect 4063 -2292 4079 -2258
rect 4137 -2292 4153 -2258
rect 4221 -2292 4237 -2258
rect 4295 -2292 4311 -2258
rect 4379 -2292 4395 -2258
rect 4453 -2292 4469 -2258
rect 4537 -2292 4553 -2258
rect 4611 -2292 4627 -2258
rect 4695 -2292 4711 -2258
rect 4769 -2292 4785 -2258
rect 4853 -2292 4869 -2258
rect 4927 -2292 4943 -2258
rect 5011 -2292 5027 -2258
rect 5085 -2292 5101 -2258
rect 5169 -2292 5185 -2258
rect 5243 -2292 5259 -2258
rect 5327 -2292 5343 -2258
rect 5401 -2292 5417 -2258
rect 5485 -2292 5501 -2258
rect 5559 -2292 5575 -2258
rect 5643 -2292 5659 -2258
rect 5717 -2292 5733 -2258
rect 5801 -2292 5817 -2258
rect 5875 -2292 5891 -2258
rect 5959 -2292 5975 -2258
rect 6033 -2292 6049 -2258
rect 6117 -2292 6133 -2258
rect 6191 -2292 6207 -2258
rect 6275 -2292 6291 -2258
rect -6471 -2396 -6437 -2334
rect 6437 -2396 6471 -2334
rect -6471 -2430 -6375 -2396
rect 6375 -2430 6471 -2396
<< viali >>
rect -6275 2258 -6207 2292
rect -6117 2258 -6049 2292
rect -5959 2258 -5891 2292
rect -5801 2258 -5733 2292
rect -5643 2258 -5575 2292
rect -5485 2258 -5417 2292
rect -5327 2258 -5259 2292
rect -5169 2258 -5101 2292
rect -5011 2258 -4943 2292
rect -4853 2258 -4785 2292
rect -4695 2258 -4627 2292
rect -4537 2258 -4469 2292
rect -4379 2258 -4311 2292
rect -4221 2258 -4153 2292
rect -4063 2258 -3995 2292
rect -3905 2258 -3837 2292
rect -3747 2258 -3679 2292
rect -3589 2258 -3521 2292
rect -3431 2258 -3363 2292
rect -3273 2258 -3205 2292
rect -3115 2258 -3047 2292
rect -2957 2258 -2889 2292
rect -2799 2258 -2731 2292
rect -2641 2258 -2573 2292
rect -2483 2258 -2415 2292
rect -2325 2258 -2257 2292
rect -2167 2258 -2099 2292
rect -2009 2258 -1941 2292
rect -1851 2258 -1783 2292
rect -1693 2258 -1625 2292
rect -1535 2258 -1467 2292
rect -1377 2258 -1309 2292
rect -1219 2258 -1151 2292
rect -1061 2258 -993 2292
rect -903 2258 -835 2292
rect -745 2258 -677 2292
rect -587 2258 -519 2292
rect -429 2258 -361 2292
rect -271 2258 -203 2292
rect -113 2258 -45 2292
rect 45 2258 113 2292
rect 203 2258 271 2292
rect 361 2258 429 2292
rect 519 2258 587 2292
rect 677 2258 745 2292
rect 835 2258 903 2292
rect 993 2258 1061 2292
rect 1151 2258 1219 2292
rect 1309 2258 1377 2292
rect 1467 2258 1535 2292
rect 1625 2258 1693 2292
rect 1783 2258 1851 2292
rect 1941 2258 2009 2292
rect 2099 2258 2167 2292
rect 2257 2258 2325 2292
rect 2415 2258 2483 2292
rect 2573 2258 2641 2292
rect 2731 2258 2799 2292
rect 2889 2258 2957 2292
rect 3047 2258 3115 2292
rect 3205 2258 3273 2292
rect 3363 2258 3431 2292
rect 3521 2258 3589 2292
rect 3679 2258 3747 2292
rect 3837 2258 3905 2292
rect 3995 2258 4063 2292
rect 4153 2258 4221 2292
rect 4311 2258 4379 2292
rect 4469 2258 4537 2292
rect 4627 2258 4695 2292
rect 4785 2258 4853 2292
rect 4943 2258 5011 2292
rect 5101 2258 5169 2292
rect 5259 2258 5327 2292
rect 5417 2258 5485 2292
rect 5575 2258 5643 2292
rect 5733 2258 5801 2292
rect 5891 2258 5959 2292
rect 6049 2258 6117 2292
rect 6207 2258 6275 2292
rect -6337 1432 -6303 2208
rect -6179 1432 -6145 2208
rect -6021 1432 -5987 2208
rect -5863 1432 -5829 2208
rect -5705 1432 -5671 2208
rect -5547 1432 -5513 2208
rect -5389 1432 -5355 2208
rect -5231 1432 -5197 2208
rect -5073 1432 -5039 2208
rect -4915 1432 -4881 2208
rect -4757 1432 -4723 2208
rect -4599 1432 -4565 2208
rect -4441 1432 -4407 2208
rect -4283 1432 -4249 2208
rect -4125 1432 -4091 2208
rect -3967 1432 -3933 2208
rect -3809 1432 -3775 2208
rect -3651 1432 -3617 2208
rect -3493 1432 -3459 2208
rect -3335 1432 -3301 2208
rect -3177 1432 -3143 2208
rect -3019 1432 -2985 2208
rect -2861 1432 -2827 2208
rect -2703 1432 -2669 2208
rect -2545 1432 -2511 2208
rect -2387 1432 -2353 2208
rect -2229 1432 -2195 2208
rect -2071 1432 -2037 2208
rect -1913 1432 -1879 2208
rect -1755 1432 -1721 2208
rect -1597 1432 -1563 2208
rect -1439 1432 -1405 2208
rect -1281 1432 -1247 2208
rect -1123 1432 -1089 2208
rect -965 1432 -931 2208
rect -807 1432 -773 2208
rect -649 1432 -615 2208
rect -491 1432 -457 2208
rect -333 1432 -299 2208
rect -175 1432 -141 2208
rect -17 1432 17 2208
rect 141 1432 175 2208
rect 299 1432 333 2208
rect 457 1432 491 2208
rect 615 1432 649 2208
rect 773 1432 807 2208
rect 931 1432 965 2208
rect 1089 1432 1123 2208
rect 1247 1432 1281 2208
rect 1405 1432 1439 2208
rect 1563 1432 1597 2208
rect 1721 1432 1755 2208
rect 1879 1432 1913 2208
rect 2037 1432 2071 2208
rect 2195 1432 2229 2208
rect 2353 1432 2387 2208
rect 2511 1432 2545 2208
rect 2669 1432 2703 2208
rect 2827 1432 2861 2208
rect 2985 1432 3019 2208
rect 3143 1432 3177 2208
rect 3301 1432 3335 2208
rect 3459 1432 3493 2208
rect 3617 1432 3651 2208
rect 3775 1432 3809 2208
rect 3933 1432 3967 2208
rect 4091 1432 4125 2208
rect 4249 1432 4283 2208
rect 4407 1432 4441 2208
rect 4565 1432 4599 2208
rect 4723 1432 4757 2208
rect 4881 1432 4915 2208
rect 5039 1432 5073 2208
rect 5197 1432 5231 2208
rect 5355 1432 5389 2208
rect 5513 1432 5547 2208
rect 5671 1432 5705 2208
rect 5829 1432 5863 2208
rect 5987 1432 6021 2208
rect 6145 1432 6179 2208
rect 6303 1432 6337 2208
rect -6275 1348 -6207 1382
rect -6117 1348 -6049 1382
rect -5959 1348 -5891 1382
rect -5801 1348 -5733 1382
rect -5643 1348 -5575 1382
rect -5485 1348 -5417 1382
rect -5327 1348 -5259 1382
rect -5169 1348 -5101 1382
rect -5011 1348 -4943 1382
rect -4853 1348 -4785 1382
rect -4695 1348 -4627 1382
rect -4537 1348 -4469 1382
rect -4379 1348 -4311 1382
rect -4221 1348 -4153 1382
rect -4063 1348 -3995 1382
rect -3905 1348 -3837 1382
rect -3747 1348 -3679 1382
rect -3589 1348 -3521 1382
rect -3431 1348 -3363 1382
rect -3273 1348 -3205 1382
rect -3115 1348 -3047 1382
rect -2957 1348 -2889 1382
rect -2799 1348 -2731 1382
rect -2641 1348 -2573 1382
rect -2483 1348 -2415 1382
rect -2325 1348 -2257 1382
rect -2167 1348 -2099 1382
rect -2009 1348 -1941 1382
rect -1851 1348 -1783 1382
rect -1693 1348 -1625 1382
rect -1535 1348 -1467 1382
rect -1377 1348 -1309 1382
rect -1219 1348 -1151 1382
rect -1061 1348 -993 1382
rect -903 1348 -835 1382
rect -745 1348 -677 1382
rect -587 1348 -519 1382
rect -429 1348 -361 1382
rect -271 1348 -203 1382
rect -113 1348 -45 1382
rect 45 1348 113 1382
rect 203 1348 271 1382
rect 361 1348 429 1382
rect 519 1348 587 1382
rect 677 1348 745 1382
rect 835 1348 903 1382
rect 993 1348 1061 1382
rect 1151 1348 1219 1382
rect 1309 1348 1377 1382
rect 1467 1348 1535 1382
rect 1625 1348 1693 1382
rect 1783 1348 1851 1382
rect 1941 1348 2009 1382
rect 2099 1348 2167 1382
rect 2257 1348 2325 1382
rect 2415 1348 2483 1382
rect 2573 1348 2641 1382
rect 2731 1348 2799 1382
rect 2889 1348 2957 1382
rect 3047 1348 3115 1382
rect 3205 1348 3273 1382
rect 3363 1348 3431 1382
rect 3521 1348 3589 1382
rect 3679 1348 3747 1382
rect 3837 1348 3905 1382
rect 3995 1348 4063 1382
rect 4153 1348 4221 1382
rect 4311 1348 4379 1382
rect 4469 1348 4537 1382
rect 4627 1348 4695 1382
rect 4785 1348 4853 1382
rect 4943 1348 5011 1382
rect 5101 1348 5169 1382
rect 5259 1348 5327 1382
rect 5417 1348 5485 1382
rect 5575 1348 5643 1382
rect 5733 1348 5801 1382
rect 5891 1348 5959 1382
rect 6049 1348 6117 1382
rect 6207 1348 6275 1382
rect -6337 522 -6303 1298
rect -6179 522 -6145 1298
rect -6021 522 -5987 1298
rect -5863 522 -5829 1298
rect -5705 522 -5671 1298
rect -5547 522 -5513 1298
rect -5389 522 -5355 1298
rect -5231 522 -5197 1298
rect -5073 522 -5039 1298
rect -4915 522 -4881 1298
rect -4757 522 -4723 1298
rect -4599 522 -4565 1298
rect -4441 522 -4407 1298
rect -4283 522 -4249 1298
rect -4125 522 -4091 1298
rect -3967 522 -3933 1298
rect -3809 522 -3775 1298
rect -3651 522 -3617 1298
rect -3493 522 -3459 1298
rect -3335 522 -3301 1298
rect -3177 522 -3143 1298
rect -3019 522 -2985 1298
rect -2861 522 -2827 1298
rect -2703 522 -2669 1298
rect -2545 522 -2511 1298
rect -2387 522 -2353 1298
rect -2229 522 -2195 1298
rect -2071 522 -2037 1298
rect -1913 522 -1879 1298
rect -1755 522 -1721 1298
rect -1597 522 -1563 1298
rect -1439 522 -1405 1298
rect -1281 522 -1247 1298
rect -1123 522 -1089 1298
rect -965 522 -931 1298
rect -807 522 -773 1298
rect -649 522 -615 1298
rect -491 522 -457 1298
rect -333 522 -299 1298
rect -175 522 -141 1298
rect -17 522 17 1298
rect 141 522 175 1298
rect 299 522 333 1298
rect 457 522 491 1298
rect 615 522 649 1298
rect 773 522 807 1298
rect 931 522 965 1298
rect 1089 522 1123 1298
rect 1247 522 1281 1298
rect 1405 522 1439 1298
rect 1563 522 1597 1298
rect 1721 522 1755 1298
rect 1879 522 1913 1298
rect 2037 522 2071 1298
rect 2195 522 2229 1298
rect 2353 522 2387 1298
rect 2511 522 2545 1298
rect 2669 522 2703 1298
rect 2827 522 2861 1298
rect 2985 522 3019 1298
rect 3143 522 3177 1298
rect 3301 522 3335 1298
rect 3459 522 3493 1298
rect 3617 522 3651 1298
rect 3775 522 3809 1298
rect 3933 522 3967 1298
rect 4091 522 4125 1298
rect 4249 522 4283 1298
rect 4407 522 4441 1298
rect 4565 522 4599 1298
rect 4723 522 4757 1298
rect 4881 522 4915 1298
rect 5039 522 5073 1298
rect 5197 522 5231 1298
rect 5355 522 5389 1298
rect 5513 522 5547 1298
rect 5671 522 5705 1298
rect 5829 522 5863 1298
rect 5987 522 6021 1298
rect 6145 522 6179 1298
rect 6303 522 6337 1298
rect -6275 438 -6207 472
rect -6117 438 -6049 472
rect -5959 438 -5891 472
rect -5801 438 -5733 472
rect -5643 438 -5575 472
rect -5485 438 -5417 472
rect -5327 438 -5259 472
rect -5169 438 -5101 472
rect -5011 438 -4943 472
rect -4853 438 -4785 472
rect -4695 438 -4627 472
rect -4537 438 -4469 472
rect -4379 438 -4311 472
rect -4221 438 -4153 472
rect -4063 438 -3995 472
rect -3905 438 -3837 472
rect -3747 438 -3679 472
rect -3589 438 -3521 472
rect -3431 438 -3363 472
rect -3273 438 -3205 472
rect -3115 438 -3047 472
rect -2957 438 -2889 472
rect -2799 438 -2731 472
rect -2641 438 -2573 472
rect -2483 438 -2415 472
rect -2325 438 -2257 472
rect -2167 438 -2099 472
rect -2009 438 -1941 472
rect -1851 438 -1783 472
rect -1693 438 -1625 472
rect -1535 438 -1467 472
rect -1377 438 -1309 472
rect -1219 438 -1151 472
rect -1061 438 -993 472
rect -903 438 -835 472
rect -745 438 -677 472
rect -587 438 -519 472
rect -429 438 -361 472
rect -271 438 -203 472
rect -113 438 -45 472
rect 45 438 113 472
rect 203 438 271 472
rect 361 438 429 472
rect 519 438 587 472
rect 677 438 745 472
rect 835 438 903 472
rect 993 438 1061 472
rect 1151 438 1219 472
rect 1309 438 1377 472
rect 1467 438 1535 472
rect 1625 438 1693 472
rect 1783 438 1851 472
rect 1941 438 2009 472
rect 2099 438 2167 472
rect 2257 438 2325 472
rect 2415 438 2483 472
rect 2573 438 2641 472
rect 2731 438 2799 472
rect 2889 438 2957 472
rect 3047 438 3115 472
rect 3205 438 3273 472
rect 3363 438 3431 472
rect 3521 438 3589 472
rect 3679 438 3747 472
rect 3837 438 3905 472
rect 3995 438 4063 472
rect 4153 438 4221 472
rect 4311 438 4379 472
rect 4469 438 4537 472
rect 4627 438 4695 472
rect 4785 438 4853 472
rect 4943 438 5011 472
rect 5101 438 5169 472
rect 5259 438 5327 472
rect 5417 438 5485 472
rect 5575 438 5643 472
rect 5733 438 5801 472
rect 5891 438 5959 472
rect 6049 438 6117 472
rect 6207 438 6275 472
rect -6337 -388 -6303 388
rect -6179 -388 -6145 388
rect -6021 -388 -5987 388
rect -5863 -388 -5829 388
rect -5705 -388 -5671 388
rect -5547 -388 -5513 388
rect -5389 -388 -5355 388
rect -5231 -388 -5197 388
rect -5073 -388 -5039 388
rect -4915 -388 -4881 388
rect -4757 -388 -4723 388
rect -4599 -388 -4565 388
rect -4441 -388 -4407 388
rect -4283 -388 -4249 388
rect -4125 -388 -4091 388
rect -3967 -388 -3933 388
rect -3809 -388 -3775 388
rect -3651 -388 -3617 388
rect -3493 -388 -3459 388
rect -3335 -388 -3301 388
rect -3177 -388 -3143 388
rect -3019 -388 -2985 388
rect -2861 -388 -2827 388
rect -2703 -388 -2669 388
rect -2545 -388 -2511 388
rect -2387 -388 -2353 388
rect -2229 -388 -2195 388
rect -2071 -388 -2037 388
rect -1913 -388 -1879 388
rect -1755 -388 -1721 388
rect -1597 -388 -1563 388
rect -1439 -388 -1405 388
rect -1281 -388 -1247 388
rect -1123 -388 -1089 388
rect -965 -388 -931 388
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
rect 931 -388 965 388
rect 1089 -388 1123 388
rect 1247 -388 1281 388
rect 1405 -388 1439 388
rect 1563 -388 1597 388
rect 1721 -388 1755 388
rect 1879 -388 1913 388
rect 2037 -388 2071 388
rect 2195 -388 2229 388
rect 2353 -388 2387 388
rect 2511 -388 2545 388
rect 2669 -388 2703 388
rect 2827 -388 2861 388
rect 2985 -388 3019 388
rect 3143 -388 3177 388
rect 3301 -388 3335 388
rect 3459 -388 3493 388
rect 3617 -388 3651 388
rect 3775 -388 3809 388
rect 3933 -388 3967 388
rect 4091 -388 4125 388
rect 4249 -388 4283 388
rect 4407 -388 4441 388
rect 4565 -388 4599 388
rect 4723 -388 4757 388
rect 4881 -388 4915 388
rect 5039 -388 5073 388
rect 5197 -388 5231 388
rect 5355 -388 5389 388
rect 5513 -388 5547 388
rect 5671 -388 5705 388
rect 5829 -388 5863 388
rect 5987 -388 6021 388
rect 6145 -388 6179 388
rect 6303 -388 6337 388
rect -6275 -472 -6207 -438
rect -6117 -472 -6049 -438
rect -5959 -472 -5891 -438
rect -5801 -472 -5733 -438
rect -5643 -472 -5575 -438
rect -5485 -472 -5417 -438
rect -5327 -472 -5259 -438
rect -5169 -472 -5101 -438
rect -5011 -472 -4943 -438
rect -4853 -472 -4785 -438
rect -4695 -472 -4627 -438
rect -4537 -472 -4469 -438
rect -4379 -472 -4311 -438
rect -4221 -472 -4153 -438
rect -4063 -472 -3995 -438
rect -3905 -472 -3837 -438
rect -3747 -472 -3679 -438
rect -3589 -472 -3521 -438
rect -3431 -472 -3363 -438
rect -3273 -472 -3205 -438
rect -3115 -472 -3047 -438
rect -2957 -472 -2889 -438
rect -2799 -472 -2731 -438
rect -2641 -472 -2573 -438
rect -2483 -472 -2415 -438
rect -2325 -472 -2257 -438
rect -2167 -472 -2099 -438
rect -2009 -472 -1941 -438
rect -1851 -472 -1783 -438
rect -1693 -472 -1625 -438
rect -1535 -472 -1467 -438
rect -1377 -472 -1309 -438
rect -1219 -472 -1151 -438
rect -1061 -472 -993 -438
rect -903 -472 -835 -438
rect -745 -472 -677 -438
rect -587 -472 -519 -438
rect -429 -472 -361 -438
rect -271 -472 -203 -438
rect -113 -472 -45 -438
rect 45 -472 113 -438
rect 203 -472 271 -438
rect 361 -472 429 -438
rect 519 -472 587 -438
rect 677 -472 745 -438
rect 835 -472 903 -438
rect 993 -472 1061 -438
rect 1151 -472 1219 -438
rect 1309 -472 1377 -438
rect 1467 -472 1535 -438
rect 1625 -472 1693 -438
rect 1783 -472 1851 -438
rect 1941 -472 2009 -438
rect 2099 -472 2167 -438
rect 2257 -472 2325 -438
rect 2415 -472 2483 -438
rect 2573 -472 2641 -438
rect 2731 -472 2799 -438
rect 2889 -472 2957 -438
rect 3047 -472 3115 -438
rect 3205 -472 3273 -438
rect 3363 -472 3431 -438
rect 3521 -472 3589 -438
rect 3679 -472 3747 -438
rect 3837 -472 3905 -438
rect 3995 -472 4063 -438
rect 4153 -472 4221 -438
rect 4311 -472 4379 -438
rect 4469 -472 4537 -438
rect 4627 -472 4695 -438
rect 4785 -472 4853 -438
rect 4943 -472 5011 -438
rect 5101 -472 5169 -438
rect 5259 -472 5327 -438
rect 5417 -472 5485 -438
rect 5575 -472 5643 -438
rect 5733 -472 5801 -438
rect 5891 -472 5959 -438
rect 6049 -472 6117 -438
rect 6207 -472 6275 -438
rect -6337 -1298 -6303 -522
rect -6179 -1298 -6145 -522
rect -6021 -1298 -5987 -522
rect -5863 -1298 -5829 -522
rect -5705 -1298 -5671 -522
rect -5547 -1298 -5513 -522
rect -5389 -1298 -5355 -522
rect -5231 -1298 -5197 -522
rect -5073 -1298 -5039 -522
rect -4915 -1298 -4881 -522
rect -4757 -1298 -4723 -522
rect -4599 -1298 -4565 -522
rect -4441 -1298 -4407 -522
rect -4283 -1298 -4249 -522
rect -4125 -1298 -4091 -522
rect -3967 -1298 -3933 -522
rect -3809 -1298 -3775 -522
rect -3651 -1298 -3617 -522
rect -3493 -1298 -3459 -522
rect -3335 -1298 -3301 -522
rect -3177 -1298 -3143 -522
rect -3019 -1298 -2985 -522
rect -2861 -1298 -2827 -522
rect -2703 -1298 -2669 -522
rect -2545 -1298 -2511 -522
rect -2387 -1298 -2353 -522
rect -2229 -1298 -2195 -522
rect -2071 -1298 -2037 -522
rect -1913 -1298 -1879 -522
rect -1755 -1298 -1721 -522
rect -1597 -1298 -1563 -522
rect -1439 -1298 -1405 -522
rect -1281 -1298 -1247 -522
rect -1123 -1298 -1089 -522
rect -965 -1298 -931 -522
rect -807 -1298 -773 -522
rect -649 -1298 -615 -522
rect -491 -1298 -457 -522
rect -333 -1298 -299 -522
rect -175 -1298 -141 -522
rect -17 -1298 17 -522
rect 141 -1298 175 -522
rect 299 -1298 333 -522
rect 457 -1298 491 -522
rect 615 -1298 649 -522
rect 773 -1298 807 -522
rect 931 -1298 965 -522
rect 1089 -1298 1123 -522
rect 1247 -1298 1281 -522
rect 1405 -1298 1439 -522
rect 1563 -1298 1597 -522
rect 1721 -1298 1755 -522
rect 1879 -1298 1913 -522
rect 2037 -1298 2071 -522
rect 2195 -1298 2229 -522
rect 2353 -1298 2387 -522
rect 2511 -1298 2545 -522
rect 2669 -1298 2703 -522
rect 2827 -1298 2861 -522
rect 2985 -1298 3019 -522
rect 3143 -1298 3177 -522
rect 3301 -1298 3335 -522
rect 3459 -1298 3493 -522
rect 3617 -1298 3651 -522
rect 3775 -1298 3809 -522
rect 3933 -1298 3967 -522
rect 4091 -1298 4125 -522
rect 4249 -1298 4283 -522
rect 4407 -1298 4441 -522
rect 4565 -1298 4599 -522
rect 4723 -1298 4757 -522
rect 4881 -1298 4915 -522
rect 5039 -1298 5073 -522
rect 5197 -1298 5231 -522
rect 5355 -1298 5389 -522
rect 5513 -1298 5547 -522
rect 5671 -1298 5705 -522
rect 5829 -1298 5863 -522
rect 5987 -1298 6021 -522
rect 6145 -1298 6179 -522
rect 6303 -1298 6337 -522
rect -6275 -1382 -6207 -1348
rect -6117 -1382 -6049 -1348
rect -5959 -1382 -5891 -1348
rect -5801 -1382 -5733 -1348
rect -5643 -1382 -5575 -1348
rect -5485 -1382 -5417 -1348
rect -5327 -1382 -5259 -1348
rect -5169 -1382 -5101 -1348
rect -5011 -1382 -4943 -1348
rect -4853 -1382 -4785 -1348
rect -4695 -1382 -4627 -1348
rect -4537 -1382 -4469 -1348
rect -4379 -1382 -4311 -1348
rect -4221 -1382 -4153 -1348
rect -4063 -1382 -3995 -1348
rect -3905 -1382 -3837 -1348
rect -3747 -1382 -3679 -1348
rect -3589 -1382 -3521 -1348
rect -3431 -1382 -3363 -1348
rect -3273 -1382 -3205 -1348
rect -3115 -1382 -3047 -1348
rect -2957 -1382 -2889 -1348
rect -2799 -1382 -2731 -1348
rect -2641 -1382 -2573 -1348
rect -2483 -1382 -2415 -1348
rect -2325 -1382 -2257 -1348
rect -2167 -1382 -2099 -1348
rect -2009 -1382 -1941 -1348
rect -1851 -1382 -1783 -1348
rect -1693 -1382 -1625 -1348
rect -1535 -1382 -1467 -1348
rect -1377 -1382 -1309 -1348
rect -1219 -1382 -1151 -1348
rect -1061 -1382 -993 -1348
rect -903 -1382 -835 -1348
rect -745 -1382 -677 -1348
rect -587 -1382 -519 -1348
rect -429 -1382 -361 -1348
rect -271 -1382 -203 -1348
rect -113 -1382 -45 -1348
rect 45 -1382 113 -1348
rect 203 -1382 271 -1348
rect 361 -1382 429 -1348
rect 519 -1382 587 -1348
rect 677 -1382 745 -1348
rect 835 -1382 903 -1348
rect 993 -1382 1061 -1348
rect 1151 -1382 1219 -1348
rect 1309 -1382 1377 -1348
rect 1467 -1382 1535 -1348
rect 1625 -1382 1693 -1348
rect 1783 -1382 1851 -1348
rect 1941 -1382 2009 -1348
rect 2099 -1382 2167 -1348
rect 2257 -1382 2325 -1348
rect 2415 -1382 2483 -1348
rect 2573 -1382 2641 -1348
rect 2731 -1382 2799 -1348
rect 2889 -1382 2957 -1348
rect 3047 -1382 3115 -1348
rect 3205 -1382 3273 -1348
rect 3363 -1382 3431 -1348
rect 3521 -1382 3589 -1348
rect 3679 -1382 3747 -1348
rect 3837 -1382 3905 -1348
rect 3995 -1382 4063 -1348
rect 4153 -1382 4221 -1348
rect 4311 -1382 4379 -1348
rect 4469 -1382 4537 -1348
rect 4627 -1382 4695 -1348
rect 4785 -1382 4853 -1348
rect 4943 -1382 5011 -1348
rect 5101 -1382 5169 -1348
rect 5259 -1382 5327 -1348
rect 5417 -1382 5485 -1348
rect 5575 -1382 5643 -1348
rect 5733 -1382 5801 -1348
rect 5891 -1382 5959 -1348
rect 6049 -1382 6117 -1348
rect 6207 -1382 6275 -1348
rect -6337 -2208 -6303 -1432
rect -6179 -2208 -6145 -1432
rect -6021 -2208 -5987 -1432
rect -5863 -2208 -5829 -1432
rect -5705 -2208 -5671 -1432
rect -5547 -2208 -5513 -1432
rect -5389 -2208 -5355 -1432
rect -5231 -2208 -5197 -1432
rect -5073 -2208 -5039 -1432
rect -4915 -2208 -4881 -1432
rect -4757 -2208 -4723 -1432
rect -4599 -2208 -4565 -1432
rect -4441 -2208 -4407 -1432
rect -4283 -2208 -4249 -1432
rect -4125 -2208 -4091 -1432
rect -3967 -2208 -3933 -1432
rect -3809 -2208 -3775 -1432
rect -3651 -2208 -3617 -1432
rect -3493 -2208 -3459 -1432
rect -3335 -2208 -3301 -1432
rect -3177 -2208 -3143 -1432
rect -3019 -2208 -2985 -1432
rect -2861 -2208 -2827 -1432
rect -2703 -2208 -2669 -1432
rect -2545 -2208 -2511 -1432
rect -2387 -2208 -2353 -1432
rect -2229 -2208 -2195 -1432
rect -2071 -2208 -2037 -1432
rect -1913 -2208 -1879 -1432
rect -1755 -2208 -1721 -1432
rect -1597 -2208 -1563 -1432
rect -1439 -2208 -1405 -1432
rect -1281 -2208 -1247 -1432
rect -1123 -2208 -1089 -1432
rect -965 -2208 -931 -1432
rect -807 -2208 -773 -1432
rect -649 -2208 -615 -1432
rect -491 -2208 -457 -1432
rect -333 -2208 -299 -1432
rect -175 -2208 -141 -1432
rect -17 -2208 17 -1432
rect 141 -2208 175 -1432
rect 299 -2208 333 -1432
rect 457 -2208 491 -1432
rect 615 -2208 649 -1432
rect 773 -2208 807 -1432
rect 931 -2208 965 -1432
rect 1089 -2208 1123 -1432
rect 1247 -2208 1281 -1432
rect 1405 -2208 1439 -1432
rect 1563 -2208 1597 -1432
rect 1721 -2208 1755 -1432
rect 1879 -2208 1913 -1432
rect 2037 -2208 2071 -1432
rect 2195 -2208 2229 -1432
rect 2353 -2208 2387 -1432
rect 2511 -2208 2545 -1432
rect 2669 -2208 2703 -1432
rect 2827 -2208 2861 -1432
rect 2985 -2208 3019 -1432
rect 3143 -2208 3177 -1432
rect 3301 -2208 3335 -1432
rect 3459 -2208 3493 -1432
rect 3617 -2208 3651 -1432
rect 3775 -2208 3809 -1432
rect 3933 -2208 3967 -1432
rect 4091 -2208 4125 -1432
rect 4249 -2208 4283 -1432
rect 4407 -2208 4441 -1432
rect 4565 -2208 4599 -1432
rect 4723 -2208 4757 -1432
rect 4881 -2208 4915 -1432
rect 5039 -2208 5073 -1432
rect 5197 -2208 5231 -1432
rect 5355 -2208 5389 -1432
rect 5513 -2208 5547 -1432
rect 5671 -2208 5705 -1432
rect 5829 -2208 5863 -1432
rect 5987 -2208 6021 -1432
rect 6145 -2208 6179 -1432
rect 6303 -2208 6337 -1432
rect -6275 -2292 -6207 -2258
rect -6117 -2292 -6049 -2258
rect -5959 -2292 -5891 -2258
rect -5801 -2292 -5733 -2258
rect -5643 -2292 -5575 -2258
rect -5485 -2292 -5417 -2258
rect -5327 -2292 -5259 -2258
rect -5169 -2292 -5101 -2258
rect -5011 -2292 -4943 -2258
rect -4853 -2292 -4785 -2258
rect -4695 -2292 -4627 -2258
rect -4537 -2292 -4469 -2258
rect -4379 -2292 -4311 -2258
rect -4221 -2292 -4153 -2258
rect -4063 -2292 -3995 -2258
rect -3905 -2292 -3837 -2258
rect -3747 -2292 -3679 -2258
rect -3589 -2292 -3521 -2258
rect -3431 -2292 -3363 -2258
rect -3273 -2292 -3205 -2258
rect -3115 -2292 -3047 -2258
rect -2957 -2292 -2889 -2258
rect -2799 -2292 -2731 -2258
rect -2641 -2292 -2573 -2258
rect -2483 -2292 -2415 -2258
rect -2325 -2292 -2257 -2258
rect -2167 -2292 -2099 -2258
rect -2009 -2292 -1941 -2258
rect -1851 -2292 -1783 -2258
rect -1693 -2292 -1625 -2258
rect -1535 -2292 -1467 -2258
rect -1377 -2292 -1309 -2258
rect -1219 -2292 -1151 -2258
rect -1061 -2292 -993 -2258
rect -903 -2292 -835 -2258
rect -745 -2292 -677 -2258
rect -587 -2292 -519 -2258
rect -429 -2292 -361 -2258
rect -271 -2292 -203 -2258
rect -113 -2292 -45 -2258
rect 45 -2292 113 -2258
rect 203 -2292 271 -2258
rect 361 -2292 429 -2258
rect 519 -2292 587 -2258
rect 677 -2292 745 -2258
rect 835 -2292 903 -2258
rect 993 -2292 1061 -2258
rect 1151 -2292 1219 -2258
rect 1309 -2292 1377 -2258
rect 1467 -2292 1535 -2258
rect 1625 -2292 1693 -2258
rect 1783 -2292 1851 -2258
rect 1941 -2292 2009 -2258
rect 2099 -2292 2167 -2258
rect 2257 -2292 2325 -2258
rect 2415 -2292 2483 -2258
rect 2573 -2292 2641 -2258
rect 2731 -2292 2799 -2258
rect 2889 -2292 2957 -2258
rect 3047 -2292 3115 -2258
rect 3205 -2292 3273 -2258
rect 3363 -2292 3431 -2258
rect 3521 -2292 3589 -2258
rect 3679 -2292 3747 -2258
rect 3837 -2292 3905 -2258
rect 3995 -2292 4063 -2258
rect 4153 -2292 4221 -2258
rect 4311 -2292 4379 -2258
rect 4469 -2292 4537 -2258
rect 4627 -2292 4695 -2258
rect 4785 -2292 4853 -2258
rect 4943 -2292 5011 -2258
rect 5101 -2292 5169 -2258
rect 5259 -2292 5327 -2258
rect 5417 -2292 5485 -2258
rect 5575 -2292 5643 -2258
rect 5733 -2292 5801 -2258
rect 5891 -2292 5959 -2258
rect 6049 -2292 6117 -2258
rect 6207 -2292 6275 -2258
<< metal1 >>
rect -6287 2292 -6195 2298
rect -6287 2258 -6275 2292
rect -6207 2258 -6195 2292
rect -6287 2252 -6195 2258
rect -6129 2292 -6037 2298
rect -6129 2258 -6117 2292
rect -6049 2258 -6037 2292
rect -6129 2252 -6037 2258
rect -5971 2292 -5879 2298
rect -5971 2258 -5959 2292
rect -5891 2258 -5879 2292
rect -5971 2252 -5879 2258
rect -5813 2292 -5721 2298
rect -5813 2258 -5801 2292
rect -5733 2258 -5721 2292
rect -5813 2252 -5721 2258
rect -5655 2292 -5563 2298
rect -5655 2258 -5643 2292
rect -5575 2258 -5563 2292
rect -5655 2252 -5563 2258
rect -5497 2292 -5405 2298
rect -5497 2258 -5485 2292
rect -5417 2258 -5405 2292
rect -5497 2252 -5405 2258
rect -5339 2292 -5247 2298
rect -5339 2258 -5327 2292
rect -5259 2258 -5247 2292
rect -5339 2252 -5247 2258
rect -5181 2292 -5089 2298
rect -5181 2258 -5169 2292
rect -5101 2258 -5089 2292
rect -5181 2252 -5089 2258
rect -5023 2292 -4931 2298
rect -5023 2258 -5011 2292
rect -4943 2258 -4931 2292
rect -5023 2252 -4931 2258
rect -4865 2292 -4773 2298
rect -4865 2258 -4853 2292
rect -4785 2258 -4773 2292
rect -4865 2252 -4773 2258
rect -4707 2292 -4615 2298
rect -4707 2258 -4695 2292
rect -4627 2258 -4615 2292
rect -4707 2252 -4615 2258
rect -4549 2292 -4457 2298
rect -4549 2258 -4537 2292
rect -4469 2258 -4457 2292
rect -4549 2252 -4457 2258
rect -4391 2292 -4299 2298
rect -4391 2258 -4379 2292
rect -4311 2258 -4299 2292
rect -4391 2252 -4299 2258
rect -4233 2292 -4141 2298
rect -4233 2258 -4221 2292
rect -4153 2258 -4141 2292
rect -4233 2252 -4141 2258
rect -4075 2292 -3983 2298
rect -4075 2258 -4063 2292
rect -3995 2258 -3983 2292
rect -4075 2252 -3983 2258
rect -3917 2292 -3825 2298
rect -3917 2258 -3905 2292
rect -3837 2258 -3825 2292
rect -3917 2252 -3825 2258
rect -3759 2292 -3667 2298
rect -3759 2258 -3747 2292
rect -3679 2258 -3667 2292
rect -3759 2252 -3667 2258
rect -3601 2292 -3509 2298
rect -3601 2258 -3589 2292
rect -3521 2258 -3509 2292
rect -3601 2252 -3509 2258
rect -3443 2292 -3351 2298
rect -3443 2258 -3431 2292
rect -3363 2258 -3351 2292
rect -3443 2252 -3351 2258
rect -3285 2292 -3193 2298
rect -3285 2258 -3273 2292
rect -3205 2258 -3193 2292
rect -3285 2252 -3193 2258
rect -3127 2292 -3035 2298
rect -3127 2258 -3115 2292
rect -3047 2258 -3035 2292
rect -3127 2252 -3035 2258
rect -2969 2292 -2877 2298
rect -2969 2258 -2957 2292
rect -2889 2258 -2877 2292
rect -2969 2252 -2877 2258
rect -2811 2292 -2719 2298
rect -2811 2258 -2799 2292
rect -2731 2258 -2719 2292
rect -2811 2252 -2719 2258
rect -2653 2292 -2561 2298
rect -2653 2258 -2641 2292
rect -2573 2258 -2561 2292
rect -2653 2252 -2561 2258
rect -2495 2292 -2403 2298
rect -2495 2258 -2483 2292
rect -2415 2258 -2403 2292
rect -2495 2252 -2403 2258
rect -2337 2292 -2245 2298
rect -2337 2258 -2325 2292
rect -2257 2258 -2245 2292
rect -2337 2252 -2245 2258
rect -2179 2292 -2087 2298
rect -2179 2258 -2167 2292
rect -2099 2258 -2087 2292
rect -2179 2252 -2087 2258
rect -2021 2292 -1929 2298
rect -2021 2258 -2009 2292
rect -1941 2258 -1929 2292
rect -2021 2252 -1929 2258
rect -1863 2292 -1771 2298
rect -1863 2258 -1851 2292
rect -1783 2258 -1771 2292
rect -1863 2252 -1771 2258
rect -1705 2292 -1613 2298
rect -1705 2258 -1693 2292
rect -1625 2258 -1613 2292
rect -1705 2252 -1613 2258
rect -1547 2292 -1455 2298
rect -1547 2258 -1535 2292
rect -1467 2258 -1455 2292
rect -1547 2252 -1455 2258
rect -1389 2292 -1297 2298
rect -1389 2258 -1377 2292
rect -1309 2258 -1297 2292
rect -1389 2252 -1297 2258
rect -1231 2292 -1139 2298
rect -1231 2258 -1219 2292
rect -1151 2258 -1139 2292
rect -1231 2252 -1139 2258
rect -1073 2292 -981 2298
rect -1073 2258 -1061 2292
rect -993 2258 -981 2292
rect -1073 2252 -981 2258
rect -915 2292 -823 2298
rect -915 2258 -903 2292
rect -835 2258 -823 2292
rect -915 2252 -823 2258
rect -757 2292 -665 2298
rect -757 2258 -745 2292
rect -677 2258 -665 2292
rect -757 2252 -665 2258
rect -599 2292 -507 2298
rect -599 2258 -587 2292
rect -519 2258 -507 2292
rect -599 2252 -507 2258
rect -441 2292 -349 2298
rect -441 2258 -429 2292
rect -361 2258 -349 2292
rect -441 2252 -349 2258
rect -283 2292 -191 2298
rect -283 2258 -271 2292
rect -203 2258 -191 2292
rect -283 2252 -191 2258
rect -125 2292 -33 2298
rect -125 2258 -113 2292
rect -45 2258 -33 2292
rect -125 2252 -33 2258
rect 33 2292 125 2298
rect 33 2258 45 2292
rect 113 2258 125 2292
rect 33 2252 125 2258
rect 191 2292 283 2298
rect 191 2258 203 2292
rect 271 2258 283 2292
rect 191 2252 283 2258
rect 349 2292 441 2298
rect 349 2258 361 2292
rect 429 2258 441 2292
rect 349 2252 441 2258
rect 507 2292 599 2298
rect 507 2258 519 2292
rect 587 2258 599 2292
rect 507 2252 599 2258
rect 665 2292 757 2298
rect 665 2258 677 2292
rect 745 2258 757 2292
rect 665 2252 757 2258
rect 823 2292 915 2298
rect 823 2258 835 2292
rect 903 2258 915 2292
rect 823 2252 915 2258
rect 981 2292 1073 2298
rect 981 2258 993 2292
rect 1061 2258 1073 2292
rect 981 2252 1073 2258
rect 1139 2292 1231 2298
rect 1139 2258 1151 2292
rect 1219 2258 1231 2292
rect 1139 2252 1231 2258
rect 1297 2292 1389 2298
rect 1297 2258 1309 2292
rect 1377 2258 1389 2292
rect 1297 2252 1389 2258
rect 1455 2292 1547 2298
rect 1455 2258 1467 2292
rect 1535 2258 1547 2292
rect 1455 2252 1547 2258
rect 1613 2292 1705 2298
rect 1613 2258 1625 2292
rect 1693 2258 1705 2292
rect 1613 2252 1705 2258
rect 1771 2292 1863 2298
rect 1771 2258 1783 2292
rect 1851 2258 1863 2292
rect 1771 2252 1863 2258
rect 1929 2292 2021 2298
rect 1929 2258 1941 2292
rect 2009 2258 2021 2292
rect 1929 2252 2021 2258
rect 2087 2292 2179 2298
rect 2087 2258 2099 2292
rect 2167 2258 2179 2292
rect 2087 2252 2179 2258
rect 2245 2292 2337 2298
rect 2245 2258 2257 2292
rect 2325 2258 2337 2292
rect 2245 2252 2337 2258
rect 2403 2292 2495 2298
rect 2403 2258 2415 2292
rect 2483 2258 2495 2292
rect 2403 2252 2495 2258
rect 2561 2292 2653 2298
rect 2561 2258 2573 2292
rect 2641 2258 2653 2292
rect 2561 2252 2653 2258
rect 2719 2292 2811 2298
rect 2719 2258 2731 2292
rect 2799 2258 2811 2292
rect 2719 2252 2811 2258
rect 2877 2292 2969 2298
rect 2877 2258 2889 2292
rect 2957 2258 2969 2292
rect 2877 2252 2969 2258
rect 3035 2292 3127 2298
rect 3035 2258 3047 2292
rect 3115 2258 3127 2292
rect 3035 2252 3127 2258
rect 3193 2292 3285 2298
rect 3193 2258 3205 2292
rect 3273 2258 3285 2292
rect 3193 2252 3285 2258
rect 3351 2292 3443 2298
rect 3351 2258 3363 2292
rect 3431 2258 3443 2292
rect 3351 2252 3443 2258
rect 3509 2292 3601 2298
rect 3509 2258 3521 2292
rect 3589 2258 3601 2292
rect 3509 2252 3601 2258
rect 3667 2292 3759 2298
rect 3667 2258 3679 2292
rect 3747 2258 3759 2292
rect 3667 2252 3759 2258
rect 3825 2292 3917 2298
rect 3825 2258 3837 2292
rect 3905 2258 3917 2292
rect 3825 2252 3917 2258
rect 3983 2292 4075 2298
rect 3983 2258 3995 2292
rect 4063 2258 4075 2292
rect 3983 2252 4075 2258
rect 4141 2292 4233 2298
rect 4141 2258 4153 2292
rect 4221 2258 4233 2292
rect 4141 2252 4233 2258
rect 4299 2292 4391 2298
rect 4299 2258 4311 2292
rect 4379 2258 4391 2292
rect 4299 2252 4391 2258
rect 4457 2292 4549 2298
rect 4457 2258 4469 2292
rect 4537 2258 4549 2292
rect 4457 2252 4549 2258
rect 4615 2292 4707 2298
rect 4615 2258 4627 2292
rect 4695 2258 4707 2292
rect 4615 2252 4707 2258
rect 4773 2292 4865 2298
rect 4773 2258 4785 2292
rect 4853 2258 4865 2292
rect 4773 2252 4865 2258
rect 4931 2292 5023 2298
rect 4931 2258 4943 2292
rect 5011 2258 5023 2292
rect 4931 2252 5023 2258
rect 5089 2292 5181 2298
rect 5089 2258 5101 2292
rect 5169 2258 5181 2292
rect 5089 2252 5181 2258
rect 5247 2292 5339 2298
rect 5247 2258 5259 2292
rect 5327 2258 5339 2292
rect 5247 2252 5339 2258
rect 5405 2292 5497 2298
rect 5405 2258 5417 2292
rect 5485 2258 5497 2292
rect 5405 2252 5497 2258
rect 5563 2292 5655 2298
rect 5563 2258 5575 2292
rect 5643 2258 5655 2292
rect 5563 2252 5655 2258
rect 5721 2292 5813 2298
rect 5721 2258 5733 2292
rect 5801 2258 5813 2292
rect 5721 2252 5813 2258
rect 5879 2292 5971 2298
rect 5879 2258 5891 2292
rect 5959 2258 5971 2292
rect 5879 2252 5971 2258
rect 6037 2292 6129 2298
rect 6037 2258 6049 2292
rect 6117 2258 6129 2292
rect 6037 2252 6129 2258
rect 6195 2292 6287 2298
rect 6195 2258 6207 2292
rect 6275 2258 6287 2292
rect 6195 2252 6287 2258
rect -6343 2208 -6297 2220
rect -6343 1432 -6337 2208
rect -6303 1432 -6297 2208
rect -6343 1420 -6297 1432
rect -6185 2208 -6139 2220
rect -6185 1432 -6179 2208
rect -6145 1432 -6139 2208
rect -6185 1420 -6139 1432
rect -6027 2208 -5981 2220
rect -6027 1432 -6021 2208
rect -5987 1432 -5981 2208
rect -6027 1420 -5981 1432
rect -5869 2208 -5823 2220
rect -5869 1432 -5863 2208
rect -5829 1432 -5823 2208
rect -5869 1420 -5823 1432
rect -5711 2208 -5665 2220
rect -5711 1432 -5705 2208
rect -5671 1432 -5665 2208
rect -5711 1420 -5665 1432
rect -5553 2208 -5507 2220
rect -5553 1432 -5547 2208
rect -5513 1432 -5507 2208
rect -5553 1420 -5507 1432
rect -5395 2208 -5349 2220
rect -5395 1432 -5389 2208
rect -5355 1432 -5349 2208
rect -5395 1420 -5349 1432
rect -5237 2208 -5191 2220
rect -5237 1432 -5231 2208
rect -5197 1432 -5191 2208
rect -5237 1420 -5191 1432
rect -5079 2208 -5033 2220
rect -5079 1432 -5073 2208
rect -5039 1432 -5033 2208
rect -5079 1420 -5033 1432
rect -4921 2208 -4875 2220
rect -4921 1432 -4915 2208
rect -4881 1432 -4875 2208
rect -4921 1420 -4875 1432
rect -4763 2208 -4717 2220
rect -4763 1432 -4757 2208
rect -4723 1432 -4717 2208
rect -4763 1420 -4717 1432
rect -4605 2208 -4559 2220
rect -4605 1432 -4599 2208
rect -4565 1432 -4559 2208
rect -4605 1420 -4559 1432
rect -4447 2208 -4401 2220
rect -4447 1432 -4441 2208
rect -4407 1432 -4401 2208
rect -4447 1420 -4401 1432
rect -4289 2208 -4243 2220
rect -4289 1432 -4283 2208
rect -4249 1432 -4243 2208
rect -4289 1420 -4243 1432
rect -4131 2208 -4085 2220
rect -4131 1432 -4125 2208
rect -4091 1432 -4085 2208
rect -4131 1420 -4085 1432
rect -3973 2208 -3927 2220
rect -3973 1432 -3967 2208
rect -3933 1432 -3927 2208
rect -3973 1420 -3927 1432
rect -3815 2208 -3769 2220
rect -3815 1432 -3809 2208
rect -3775 1432 -3769 2208
rect -3815 1420 -3769 1432
rect -3657 2208 -3611 2220
rect -3657 1432 -3651 2208
rect -3617 1432 -3611 2208
rect -3657 1420 -3611 1432
rect -3499 2208 -3453 2220
rect -3499 1432 -3493 2208
rect -3459 1432 -3453 2208
rect -3499 1420 -3453 1432
rect -3341 2208 -3295 2220
rect -3341 1432 -3335 2208
rect -3301 1432 -3295 2208
rect -3341 1420 -3295 1432
rect -3183 2208 -3137 2220
rect -3183 1432 -3177 2208
rect -3143 1432 -3137 2208
rect -3183 1420 -3137 1432
rect -3025 2208 -2979 2220
rect -3025 1432 -3019 2208
rect -2985 1432 -2979 2208
rect -3025 1420 -2979 1432
rect -2867 2208 -2821 2220
rect -2867 1432 -2861 2208
rect -2827 1432 -2821 2208
rect -2867 1420 -2821 1432
rect -2709 2208 -2663 2220
rect -2709 1432 -2703 2208
rect -2669 1432 -2663 2208
rect -2709 1420 -2663 1432
rect -2551 2208 -2505 2220
rect -2551 1432 -2545 2208
rect -2511 1432 -2505 2208
rect -2551 1420 -2505 1432
rect -2393 2208 -2347 2220
rect -2393 1432 -2387 2208
rect -2353 1432 -2347 2208
rect -2393 1420 -2347 1432
rect -2235 2208 -2189 2220
rect -2235 1432 -2229 2208
rect -2195 1432 -2189 2208
rect -2235 1420 -2189 1432
rect -2077 2208 -2031 2220
rect -2077 1432 -2071 2208
rect -2037 1432 -2031 2208
rect -2077 1420 -2031 1432
rect -1919 2208 -1873 2220
rect -1919 1432 -1913 2208
rect -1879 1432 -1873 2208
rect -1919 1420 -1873 1432
rect -1761 2208 -1715 2220
rect -1761 1432 -1755 2208
rect -1721 1432 -1715 2208
rect -1761 1420 -1715 1432
rect -1603 2208 -1557 2220
rect -1603 1432 -1597 2208
rect -1563 1432 -1557 2208
rect -1603 1420 -1557 1432
rect -1445 2208 -1399 2220
rect -1445 1432 -1439 2208
rect -1405 1432 -1399 2208
rect -1445 1420 -1399 1432
rect -1287 2208 -1241 2220
rect -1287 1432 -1281 2208
rect -1247 1432 -1241 2208
rect -1287 1420 -1241 1432
rect -1129 2208 -1083 2220
rect -1129 1432 -1123 2208
rect -1089 1432 -1083 2208
rect -1129 1420 -1083 1432
rect -971 2208 -925 2220
rect -971 1432 -965 2208
rect -931 1432 -925 2208
rect -971 1420 -925 1432
rect -813 2208 -767 2220
rect -813 1432 -807 2208
rect -773 1432 -767 2208
rect -813 1420 -767 1432
rect -655 2208 -609 2220
rect -655 1432 -649 2208
rect -615 1432 -609 2208
rect -655 1420 -609 1432
rect -497 2208 -451 2220
rect -497 1432 -491 2208
rect -457 1432 -451 2208
rect -497 1420 -451 1432
rect -339 2208 -293 2220
rect -339 1432 -333 2208
rect -299 1432 -293 2208
rect -339 1420 -293 1432
rect -181 2208 -135 2220
rect -181 1432 -175 2208
rect -141 1432 -135 2208
rect -181 1420 -135 1432
rect -23 2208 23 2220
rect -23 1432 -17 2208
rect 17 1432 23 2208
rect -23 1420 23 1432
rect 135 2208 181 2220
rect 135 1432 141 2208
rect 175 1432 181 2208
rect 135 1420 181 1432
rect 293 2208 339 2220
rect 293 1432 299 2208
rect 333 1432 339 2208
rect 293 1420 339 1432
rect 451 2208 497 2220
rect 451 1432 457 2208
rect 491 1432 497 2208
rect 451 1420 497 1432
rect 609 2208 655 2220
rect 609 1432 615 2208
rect 649 1432 655 2208
rect 609 1420 655 1432
rect 767 2208 813 2220
rect 767 1432 773 2208
rect 807 1432 813 2208
rect 767 1420 813 1432
rect 925 2208 971 2220
rect 925 1432 931 2208
rect 965 1432 971 2208
rect 925 1420 971 1432
rect 1083 2208 1129 2220
rect 1083 1432 1089 2208
rect 1123 1432 1129 2208
rect 1083 1420 1129 1432
rect 1241 2208 1287 2220
rect 1241 1432 1247 2208
rect 1281 1432 1287 2208
rect 1241 1420 1287 1432
rect 1399 2208 1445 2220
rect 1399 1432 1405 2208
rect 1439 1432 1445 2208
rect 1399 1420 1445 1432
rect 1557 2208 1603 2220
rect 1557 1432 1563 2208
rect 1597 1432 1603 2208
rect 1557 1420 1603 1432
rect 1715 2208 1761 2220
rect 1715 1432 1721 2208
rect 1755 1432 1761 2208
rect 1715 1420 1761 1432
rect 1873 2208 1919 2220
rect 1873 1432 1879 2208
rect 1913 1432 1919 2208
rect 1873 1420 1919 1432
rect 2031 2208 2077 2220
rect 2031 1432 2037 2208
rect 2071 1432 2077 2208
rect 2031 1420 2077 1432
rect 2189 2208 2235 2220
rect 2189 1432 2195 2208
rect 2229 1432 2235 2208
rect 2189 1420 2235 1432
rect 2347 2208 2393 2220
rect 2347 1432 2353 2208
rect 2387 1432 2393 2208
rect 2347 1420 2393 1432
rect 2505 2208 2551 2220
rect 2505 1432 2511 2208
rect 2545 1432 2551 2208
rect 2505 1420 2551 1432
rect 2663 2208 2709 2220
rect 2663 1432 2669 2208
rect 2703 1432 2709 2208
rect 2663 1420 2709 1432
rect 2821 2208 2867 2220
rect 2821 1432 2827 2208
rect 2861 1432 2867 2208
rect 2821 1420 2867 1432
rect 2979 2208 3025 2220
rect 2979 1432 2985 2208
rect 3019 1432 3025 2208
rect 2979 1420 3025 1432
rect 3137 2208 3183 2220
rect 3137 1432 3143 2208
rect 3177 1432 3183 2208
rect 3137 1420 3183 1432
rect 3295 2208 3341 2220
rect 3295 1432 3301 2208
rect 3335 1432 3341 2208
rect 3295 1420 3341 1432
rect 3453 2208 3499 2220
rect 3453 1432 3459 2208
rect 3493 1432 3499 2208
rect 3453 1420 3499 1432
rect 3611 2208 3657 2220
rect 3611 1432 3617 2208
rect 3651 1432 3657 2208
rect 3611 1420 3657 1432
rect 3769 2208 3815 2220
rect 3769 1432 3775 2208
rect 3809 1432 3815 2208
rect 3769 1420 3815 1432
rect 3927 2208 3973 2220
rect 3927 1432 3933 2208
rect 3967 1432 3973 2208
rect 3927 1420 3973 1432
rect 4085 2208 4131 2220
rect 4085 1432 4091 2208
rect 4125 1432 4131 2208
rect 4085 1420 4131 1432
rect 4243 2208 4289 2220
rect 4243 1432 4249 2208
rect 4283 1432 4289 2208
rect 4243 1420 4289 1432
rect 4401 2208 4447 2220
rect 4401 1432 4407 2208
rect 4441 1432 4447 2208
rect 4401 1420 4447 1432
rect 4559 2208 4605 2220
rect 4559 1432 4565 2208
rect 4599 1432 4605 2208
rect 4559 1420 4605 1432
rect 4717 2208 4763 2220
rect 4717 1432 4723 2208
rect 4757 1432 4763 2208
rect 4717 1420 4763 1432
rect 4875 2208 4921 2220
rect 4875 1432 4881 2208
rect 4915 1432 4921 2208
rect 4875 1420 4921 1432
rect 5033 2208 5079 2220
rect 5033 1432 5039 2208
rect 5073 1432 5079 2208
rect 5033 1420 5079 1432
rect 5191 2208 5237 2220
rect 5191 1432 5197 2208
rect 5231 1432 5237 2208
rect 5191 1420 5237 1432
rect 5349 2208 5395 2220
rect 5349 1432 5355 2208
rect 5389 1432 5395 2208
rect 5349 1420 5395 1432
rect 5507 2208 5553 2220
rect 5507 1432 5513 2208
rect 5547 1432 5553 2208
rect 5507 1420 5553 1432
rect 5665 2208 5711 2220
rect 5665 1432 5671 2208
rect 5705 1432 5711 2208
rect 5665 1420 5711 1432
rect 5823 2208 5869 2220
rect 5823 1432 5829 2208
rect 5863 1432 5869 2208
rect 5823 1420 5869 1432
rect 5981 2208 6027 2220
rect 5981 1432 5987 2208
rect 6021 1432 6027 2208
rect 5981 1420 6027 1432
rect 6139 2208 6185 2220
rect 6139 1432 6145 2208
rect 6179 1432 6185 2208
rect 6139 1420 6185 1432
rect 6297 2208 6343 2220
rect 6297 1432 6303 2208
rect 6337 1432 6343 2208
rect 6297 1420 6343 1432
rect -6287 1382 -6195 1388
rect -6287 1348 -6275 1382
rect -6207 1348 -6195 1382
rect -6287 1342 -6195 1348
rect -6129 1382 -6037 1388
rect -6129 1348 -6117 1382
rect -6049 1348 -6037 1382
rect -6129 1342 -6037 1348
rect -5971 1382 -5879 1388
rect -5971 1348 -5959 1382
rect -5891 1348 -5879 1382
rect -5971 1342 -5879 1348
rect -5813 1382 -5721 1388
rect -5813 1348 -5801 1382
rect -5733 1348 -5721 1382
rect -5813 1342 -5721 1348
rect -5655 1382 -5563 1388
rect -5655 1348 -5643 1382
rect -5575 1348 -5563 1382
rect -5655 1342 -5563 1348
rect -5497 1382 -5405 1388
rect -5497 1348 -5485 1382
rect -5417 1348 -5405 1382
rect -5497 1342 -5405 1348
rect -5339 1382 -5247 1388
rect -5339 1348 -5327 1382
rect -5259 1348 -5247 1382
rect -5339 1342 -5247 1348
rect -5181 1382 -5089 1388
rect -5181 1348 -5169 1382
rect -5101 1348 -5089 1382
rect -5181 1342 -5089 1348
rect -5023 1382 -4931 1388
rect -5023 1348 -5011 1382
rect -4943 1348 -4931 1382
rect -5023 1342 -4931 1348
rect -4865 1382 -4773 1388
rect -4865 1348 -4853 1382
rect -4785 1348 -4773 1382
rect -4865 1342 -4773 1348
rect -4707 1382 -4615 1388
rect -4707 1348 -4695 1382
rect -4627 1348 -4615 1382
rect -4707 1342 -4615 1348
rect -4549 1382 -4457 1388
rect -4549 1348 -4537 1382
rect -4469 1348 -4457 1382
rect -4549 1342 -4457 1348
rect -4391 1382 -4299 1388
rect -4391 1348 -4379 1382
rect -4311 1348 -4299 1382
rect -4391 1342 -4299 1348
rect -4233 1382 -4141 1388
rect -4233 1348 -4221 1382
rect -4153 1348 -4141 1382
rect -4233 1342 -4141 1348
rect -4075 1382 -3983 1388
rect -4075 1348 -4063 1382
rect -3995 1348 -3983 1382
rect -4075 1342 -3983 1348
rect -3917 1382 -3825 1388
rect -3917 1348 -3905 1382
rect -3837 1348 -3825 1382
rect -3917 1342 -3825 1348
rect -3759 1382 -3667 1388
rect -3759 1348 -3747 1382
rect -3679 1348 -3667 1382
rect -3759 1342 -3667 1348
rect -3601 1382 -3509 1388
rect -3601 1348 -3589 1382
rect -3521 1348 -3509 1382
rect -3601 1342 -3509 1348
rect -3443 1382 -3351 1388
rect -3443 1348 -3431 1382
rect -3363 1348 -3351 1382
rect -3443 1342 -3351 1348
rect -3285 1382 -3193 1388
rect -3285 1348 -3273 1382
rect -3205 1348 -3193 1382
rect -3285 1342 -3193 1348
rect -3127 1382 -3035 1388
rect -3127 1348 -3115 1382
rect -3047 1348 -3035 1382
rect -3127 1342 -3035 1348
rect -2969 1382 -2877 1388
rect -2969 1348 -2957 1382
rect -2889 1348 -2877 1382
rect -2969 1342 -2877 1348
rect -2811 1382 -2719 1388
rect -2811 1348 -2799 1382
rect -2731 1348 -2719 1382
rect -2811 1342 -2719 1348
rect -2653 1382 -2561 1388
rect -2653 1348 -2641 1382
rect -2573 1348 -2561 1382
rect -2653 1342 -2561 1348
rect -2495 1382 -2403 1388
rect -2495 1348 -2483 1382
rect -2415 1348 -2403 1382
rect -2495 1342 -2403 1348
rect -2337 1382 -2245 1388
rect -2337 1348 -2325 1382
rect -2257 1348 -2245 1382
rect -2337 1342 -2245 1348
rect -2179 1382 -2087 1388
rect -2179 1348 -2167 1382
rect -2099 1348 -2087 1382
rect -2179 1342 -2087 1348
rect -2021 1382 -1929 1388
rect -2021 1348 -2009 1382
rect -1941 1348 -1929 1382
rect -2021 1342 -1929 1348
rect -1863 1382 -1771 1388
rect -1863 1348 -1851 1382
rect -1783 1348 -1771 1382
rect -1863 1342 -1771 1348
rect -1705 1382 -1613 1388
rect -1705 1348 -1693 1382
rect -1625 1348 -1613 1382
rect -1705 1342 -1613 1348
rect -1547 1382 -1455 1388
rect -1547 1348 -1535 1382
rect -1467 1348 -1455 1382
rect -1547 1342 -1455 1348
rect -1389 1382 -1297 1388
rect -1389 1348 -1377 1382
rect -1309 1348 -1297 1382
rect -1389 1342 -1297 1348
rect -1231 1382 -1139 1388
rect -1231 1348 -1219 1382
rect -1151 1348 -1139 1382
rect -1231 1342 -1139 1348
rect -1073 1382 -981 1388
rect -1073 1348 -1061 1382
rect -993 1348 -981 1382
rect -1073 1342 -981 1348
rect -915 1382 -823 1388
rect -915 1348 -903 1382
rect -835 1348 -823 1382
rect -915 1342 -823 1348
rect -757 1382 -665 1388
rect -757 1348 -745 1382
rect -677 1348 -665 1382
rect -757 1342 -665 1348
rect -599 1382 -507 1388
rect -599 1348 -587 1382
rect -519 1348 -507 1382
rect -599 1342 -507 1348
rect -441 1382 -349 1388
rect -441 1348 -429 1382
rect -361 1348 -349 1382
rect -441 1342 -349 1348
rect -283 1382 -191 1388
rect -283 1348 -271 1382
rect -203 1348 -191 1382
rect -283 1342 -191 1348
rect -125 1382 -33 1388
rect -125 1348 -113 1382
rect -45 1348 -33 1382
rect -125 1342 -33 1348
rect 33 1382 125 1388
rect 33 1348 45 1382
rect 113 1348 125 1382
rect 33 1342 125 1348
rect 191 1382 283 1388
rect 191 1348 203 1382
rect 271 1348 283 1382
rect 191 1342 283 1348
rect 349 1382 441 1388
rect 349 1348 361 1382
rect 429 1348 441 1382
rect 349 1342 441 1348
rect 507 1382 599 1388
rect 507 1348 519 1382
rect 587 1348 599 1382
rect 507 1342 599 1348
rect 665 1382 757 1388
rect 665 1348 677 1382
rect 745 1348 757 1382
rect 665 1342 757 1348
rect 823 1382 915 1388
rect 823 1348 835 1382
rect 903 1348 915 1382
rect 823 1342 915 1348
rect 981 1382 1073 1388
rect 981 1348 993 1382
rect 1061 1348 1073 1382
rect 981 1342 1073 1348
rect 1139 1382 1231 1388
rect 1139 1348 1151 1382
rect 1219 1348 1231 1382
rect 1139 1342 1231 1348
rect 1297 1382 1389 1388
rect 1297 1348 1309 1382
rect 1377 1348 1389 1382
rect 1297 1342 1389 1348
rect 1455 1382 1547 1388
rect 1455 1348 1467 1382
rect 1535 1348 1547 1382
rect 1455 1342 1547 1348
rect 1613 1382 1705 1388
rect 1613 1348 1625 1382
rect 1693 1348 1705 1382
rect 1613 1342 1705 1348
rect 1771 1382 1863 1388
rect 1771 1348 1783 1382
rect 1851 1348 1863 1382
rect 1771 1342 1863 1348
rect 1929 1382 2021 1388
rect 1929 1348 1941 1382
rect 2009 1348 2021 1382
rect 1929 1342 2021 1348
rect 2087 1382 2179 1388
rect 2087 1348 2099 1382
rect 2167 1348 2179 1382
rect 2087 1342 2179 1348
rect 2245 1382 2337 1388
rect 2245 1348 2257 1382
rect 2325 1348 2337 1382
rect 2245 1342 2337 1348
rect 2403 1382 2495 1388
rect 2403 1348 2415 1382
rect 2483 1348 2495 1382
rect 2403 1342 2495 1348
rect 2561 1382 2653 1388
rect 2561 1348 2573 1382
rect 2641 1348 2653 1382
rect 2561 1342 2653 1348
rect 2719 1382 2811 1388
rect 2719 1348 2731 1382
rect 2799 1348 2811 1382
rect 2719 1342 2811 1348
rect 2877 1382 2969 1388
rect 2877 1348 2889 1382
rect 2957 1348 2969 1382
rect 2877 1342 2969 1348
rect 3035 1382 3127 1388
rect 3035 1348 3047 1382
rect 3115 1348 3127 1382
rect 3035 1342 3127 1348
rect 3193 1382 3285 1388
rect 3193 1348 3205 1382
rect 3273 1348 3285 1382
rect 3193 1342 3285 1348
rect 3351 1382 3443 1388
rect 3351 1348 3363 1382
rect 3431 1348 3443 1382
rect 3351 1342 3443 1348
rect 3509 1382 3601 1388
rect 3509 1348 3521 1382
rect 3589 1348 3601 1382
rect 3509 1342 3601 1348
rect 3667 1382 3759 1388
rect 3667 1348 3679 1382
rect 3747 1348 3759 1382
rect 3667 1342 3759 1348
rect 3825 1382 3917 1388
rect 3825 1348 3837 1382
rect 3905 1348 3917 1382
rect 3825 1342 3917 1348
rect 3983 1382 4075 1388
rect 3983 1348 3995 1382
rect 4063 1348 4075 1382
rect 3983 1342 4075 1348
rect 4141 1382 4233 1388
rect 4141 1348 4153 1382
rect 4221 1348 4233 1382
rect 4141 1342 4233 1348
rect 4299 1382 4391 1388
rect 4299 1348 4311 1382
rect 4379 1348 4391 1382
rect 4299 1342 4391 1348
rect 4457 1382 4549 1388
rect 4457 1348 4469 1382
rect 4537 1348 4549 1382
rect 4457 1342 4549 1348
rect 4615 1382 4707 1388
rect 4615 1348 4627 1382
rect 4695 1348 4707 1382
rect 4615 1342 4707 1348
rect 4773 1382 4865 1388
rect 4773 1348 4785 1382
rect 4853 1348 4865 1382
rect 4773 1342 4865 1348
rect 4931 1382 5023 1388
rect 4931 1348 4943 1382
rect 5011 1348 5023 1382
rect 4931 1342 5023 1348
rect 5089 1382 5181 1388
rect 5089 1348 5101 1382
rect 5169 1348 5181 1382
rect 5089 1342 5181 1348
rect 5247 1382 5339 1388
rect 5247 1348 5259 1382
rect 5327 1348 5339 1382
rect 5247 1342 5339 1348
rect 5405 1382 5497 1388
rect 5405 1348 5417 1382
rect 5485 1348 5497 1382
rect 5405 1342 5497 1348
rect 5563 1382 5655 1388
rect 5563 1348 5575 1382
rect 5643 1348 5655 1382
rect 5563 1342 5655 1348
rect 5721 1382 5813 1388
rect 5721 1348 5733 1382
rect 5801 1348 5813 1382
rect 5721 1342 5813 1348
rect 5879 1382 5971 1388
rect 5879 1348 5891 1382
rect 5959 1348 5971 1382
rect 5879 1342 5971 1348
rect 6037 1382 6129 1388
rect 6037 1348 6049 1382
rect 6117 1348 6129 1382
rect 6037 1342 6129 1348
rect 6195 1382 6287 1388
rect 6195 1348 6207 1382
rect 6275 1348 6287 1382
rect 6195 1342 6287 1348
rect -6343 1298 -6297 1310
rect -6343 522 -6337 1298
rect -6303 522 -6297 1298
rect -6343 510 -6297 522
rect -6185 1298 -6139 1310
rect -6185 522 -6179 1298
rect -6145 522 -6139 1298
rect -6185 510 -6139 522
rect -6027 1298 -5981 1310
rect -6027 522 -6021 1298
rect -5987 522 -5981 1298
rect -6027 510 -5981 522
rect -5869 1298 -5823 1310
rect -5869 522 -5863 1298
rect -5829 522 -5823 1298
rect -5869 510 -5823 522
rect -5711 1298 -5665 1310
rect -5711 522 -5705 1298
rect -5671 522 -5665 1298
rect -5711 510 -5665 522
rect -5553 1298 -5507 1310
rect -5553 522 -5547 1298
rect -5513 522 -5507 1298
rect -5553 510 -5507 522
rect -5395 1298 -5349 1310
rect -5395 522 -5389 1298
rect -5355 522 -5349 1298
rect -5395 510 -5349 522
rect -5237 1298 -5191 1310
rect -5237 522 -5231 1298
rect -5197 522 -5191 1298
rect -5237 510 -5191 522
rect -5079 1298 -5033 1310
rect -5079 522 -5073 1298
rect -5039 522 -5033 1298
rect -5079 510 -5033 522
rect -4921 1298 -4875 1310
rect -4921 522 -4915 1298
rect -4881 522 -4875 1298
rect -4921 510 -4875 522
rect -4763 1298 -4717 1310
rect -4763 522 -4757 1298
rect -4723 522 -4717 1298
rect -4763 510 -4717 522
rect -4605 1298 -4559 1310
rect -4605 522 -4599 1298
rect -4565 522 -4559 1298
rect -4605 510 -4559 522
rect -4447 1298 -4401 1310
rect -4447 522 -4441 1298
rect -4407 522 -4401 1298
rect -4447 510 -4401 522
rect -4289 1298 -4243 1310
rect -4289 522 -4283 1298
rect -4249 522 -4243 1298
rect -4289 510 -4243 522
rect -4131 1298 -4085 1310
rect -4131 522 -4125 1298
rect -4091 522 -4085 1298
rect -4131 510 -4085 522
rect -3973 1298 -3927 1310
rect -3973 522 -3967 1298
rect -3933 522 -3927 1298
rect -3973 510 -3927 522
rect -3815 1298 -3769 1310
rect -3815 522 -3809 1298
rect -3775 522 -3769 1298
rect -3815 510 -3769 522
rect -3657 1298 -3611 1310
rect -3657 522 -3651 1298
rect -3617 522 -3611 1298
rect -3657 510 -3611 522
rect -3499 1298 -3453 1310
rect -3499 522 -3493 1298
rect -3459 522 -3453 1298
rect -3499 510 -3453 522
rect -3341 1298 -3295 1310
rect -3341 522 -3335 1298
rect -3301 522 -3295 1298
rect -3341 510 -3295 522
rect -3183 1298 -3137 1310
rect -3183 522 -3177 1298
rect -3143 522 -3137 1298
rect -3183 510 -3137 522
rect -3025 1298 -2979 1310
rect -3025 522 -3019 1298
rect -2985 522 -2979 1298
rect -3025 510 -2979 522
rect -2867 1298 -2821 1310
rect -2867 522 -2861 1298
rect -2827 522 -2821 1298
rect -2867 510 -2821 522
rect -2709 1298 -2663 1310
rect -2709 522 -2703 1298
rect -2669 522 -2663 1298
rect -2709 510 -2663 522
rect -2551 1298 -2505 1310
rect -2551 522 -2545 1298
rect -2511 522 -2505 1298
rect -2551 510 -2505 522
rect -2393 1298 -2347 1310
rect -2393 522 -2387 1298
rect -2353 522 -2347 1298
rect -2393 510 -2347 522
rect -2235 1298 -2189 1310
rect -2235 522 -2229 1298
rect -2195 522 -2189 1298
rect -2235 510 -2189 522
rect -2077 1298 -2031 1310
rect -2077 522 -2071 1298
rect -2037 522 -2031 1298
rect -2077 510 -2031 522
rect -1919 1298 -1873 1310
rect -1919 522 -1913 1298
rect -1879 522 -1873 1298
rect -1919 510 -1873 522
rect -1761 1298 -1715 1310
rect -1761 522 -1755 1298
rect -1721 522 -1715 1298
rect -1761 510 -1715 522
rect -1603 1298 -1557 1310
rect -1603 522 -1597 1298
rect -1563 522 -1557 1298
rect -1603 510 -1557 522
rect -1445 1298 -1399 1310
rect -1445 522 -1439 1298
rect -1405 522 -1399 1298
rect -1445 510 -1399 522
rect -1287 1298 -1241 1310
rect -1287 522 -1281 1298
rect -1247 522 -1241 1298
rect -1287 510 -1241 522
rect -1129 1298 -1083 1310
rect -1129 522 -1123 1298
rect -1089 522 -1083 1298
rect -1129 510 -1083 522
rect -971 1298 -925 1310
rect -971 522 -965 1298
rect -931 522 -925 1298
rect -971 510 -925 522
rect -813 1298 -767 1310
rect -813 522 -807 1298
rect -773 522 -767 1298
rect -813 510 -767 522
rect -655 1298 -609 1310
rect -655 522 -649 1298
rect -615 522 -609 1298
rect -655 510 -609 522
rect -497 1298 -451 1310
rect -497 522 -491 1298
rect -457 522 -451 1298
rect -497 510 -451 522
rect -339 1298 -293 1310
rect -339 522 -333 1298
rect -299 522 -293 1298
rect -339 510 -293 522
rect -181 1298 -135 1310
rect -181 522 -175 1298
rect -141 522 -135 1298
rect -181 510 -135 522
rect -23 1298 23 1310
rect -23 522 -17 1298
rect 17 522 23 1298
rect -23 510 23 522
rect 135 1298 181 1310
rect 135 522 141 1298
rect 175 522 181 1298
rect 135 510 181 522
rect 293 1298 339 1310
rect 293 522 299 1298
rect 333 522 339 1298
rect 293 510 339 522
rect 451 1298 497 1310
rect 451 522 457 1298
rect 491 522 497 1298
rect 451 510 497 522
rect 609 1298 655 1310
rect 609 522 615 1298
rect 649 522 655 1298
rect 609 510 655 522
rect 767 1298 813 1310
rect 767 522 773 1298
rect 807 522 813 1298
rect 767 510 813 522
rect 925 1298 971 1310
rect 925 522 931 1298
rect 965 522 971 1298
rect 925 510 971 522
rect 1083 1298 1129 1310
rect 1083 522 1089 1298
rect 1123 522 1129 1298
rect 1083 510 1129 522
rect 1241 1298 1287 1310
rect 1241 522 1247 1298
rect 1281 522 1287 1298
rect 1241 510 1287 522
rect 1399 1298 1445 1310
rect 1399 522 1405 1298
rect 1439 522 1445 1298
rect 1399 510 1445 522
rect 1557 1298 1603 1310
rect 1557 522 1563 1298
rect 1597 522 1603 1298
rect 1557 510 1603 522
rect 1715 1298 1761 1310
rect 1715 522 1721 1298
rect 1755 522 1761 1298
rect 1715 510 1761 522
rect 1873 1298 1919 1310
rect 1873 522 1879 1298
rect 1913 522 1919 1298
rect 1873 510 1919 522
rect 2031 1298 2077 1310
rect 2031 522 2037 1298
rect 2071 522 2077 1298
rect 2031 510 2077 522
rect 2189 1298 2235 1310
rect 2189 522 2195 1298
rect 2229 522 2235 1298
rect 2189 510 2235 522
rect 2347 1298 2393 1310
rect 2347 522 2353 1298
rect 2387 522 2393 1298
rect 2347 510 2393 522
rect 2505 1298 2551 1310
rect 2505 522 2511 1298
rect 2545 522 2551 1298
rect 2505 510 2551 522
rect 2663 1298 2709 1310
rect 2663 522 2669 1298
rect 2703 522 2709 1298
rect 2663 510 2709 522
rect 2821 1298 2867 1310
rect 2821 522 2827 1298
rect 2861 522 2867 1298
rect 2821 510 2867 522
rect 2979 1298 3025 1310
rect 2979 522 2985 1298
rect 3019 522 3025 1298
rect 2979 510 3025 522
rect 3137 1298 3183 1310
rect 3137 522 3143 1298
rect 3177 522 3183 1298
rect 3137 510 3183 522
rect 3295 1298 3341 1310
rect 3295 522 3301 1298
rect 3335 522 3341 1298
rect 3295 510 3341 522
rect 3453 1298 3499 1310
rect 3453 522 3459 1298
rect 3493 522 3499 1298
rect 3453 510 3499 522
rect 3611 1298 3657 1310
rect 3611 522 3617 1298
rect 3651 522 3657 1298
rect 3611 510 3657 522
rect 3769 1298 3815 1310
rect 3769 522 3775 1298
rect 3809 522 3815 1298
rect 3769 510 3815 522
rect 3927 1298 3973 1310
rect 3927 522 3933 1298
rect 3967 522 3973 1298
rect 3927 510 3973 522
rect 4085 1298 4131 1310
rect 4085 522 4091 1298
rect 4125 522 4131 1298
rect 4085 510 4131 522
rect 4243 1298 4289 1310
rect 4243 522 4249 1298
rect 4283 522 4289 1298
rect 4243 510 4289 522
rect 4401 1298 4447 1310
rect 4401 522 4407 1298
rect 4441 522 4447 1298
rect 4401 510 4447 522
rect 4559 1298 4605 1310
rect 4559 522 4565 1298
rect 4599 522 4605 1298
rect 4559 510 4605 522
rect 4717 1298 4763 1310
rect 4717 522 4723 1298
rect 4757 522 4763 1298
rect 4717 510 4763 522
rect 4875 1298 4921 1310
rect 4875 522 4881 1298
rect 4915 522 4921 1298
rect 4875 510 4921 522
rect 5033 1298 5079 1310
rect 5033 522 5039 1298
rect 5073 522 5079 1298
rect 5033 510 5079 522
rect 5191 1298 5237 1310
rect 5191 522 5197 1298
rect 5231 522 5237 1298
rect 5191 510 5237 522
rect 5349 1298 5395 1310
rect 5349 522 5355 1298
rect 5389 522 5395 1298
rect 5349 510 5395 522
rect 5507 1298 5553 1310
rect 5507 522 5513 1298
rect 5547 522 5553 1298
rect 5507 510 5553 522
rect 5665 1298 5711 1310
rect 5665 522 5671 1298
rect 5705 522 5711 1298
rect 5665 510 5711 522
rect 5823 1298 5869 1310
rect 5823 522 5829 1298
rect 5863 522 5869 1298
rect 5823 510 5869 522
rect 5981 1298 6027 1310
rect 5981 522 5987 1298
rect 6021 522 6027 1298
rect 5981 510 6027 522
rect 6139 1298 6185 1310
rect 6139 522 6145 1298
rect 6179 522 6185 1298
rect 6139 510 6185 522
rect 6297 1298 6343 1310
rect 6297 522 6303 1298
rect 6337 522 6343 1298
rect 6297 510 6343 522
rect -6287 472 -6195 478
rect -6287 438 -6275 472
rect -6207 438 -6195 472
rect -6287 432 -6195 438
rect -6129 472 -6037 478
rect -6129 438 -6117 472
rect -6049 438 -6037 472
rect -6129 432 -6037 438
rect -5971 472 -5879 478
rect -5971 438 -5959 472
rect -5891 438 -5879 472
rect -5971 432 -5879 438
rect -5813 472 -5721 478
rect -5813 438 -5801 472
rect -5733 438 -5721 472
rect -5813 432 -5721 438
rect -5655 472 -5563 478
rect -5655 438 -5643 472
rect -5575 438 -5563 472
rect -5655 432 -5563 438
rect -5497 472 -5405 478
rect -5497 438 -5485 472
rect -5417 438 -5405 472
rect -5497 432 -5405 438
rect -5339 472 -5247 478
rect -5339 438 -5327 472
rect -5259 438 -5247 472
rect -5339 432 -5247 438
rect -5181 472 -5089 478
rect -5181 438 -5169 472
rect -5101 438 -5089 472
rect -5181 432 -5089 438
rect -5023 472 -4931 478
rect -5023 438 -5011 472
rect -4943 438 -4931 472
rect -5023 432 -4931 438
rect -4865 472 -4773 478
rect -4865 438 -4853 472
rect -4785 438 -4773 472
rect -4865 432 -4773 438
rect -4707 472 -4615 478
rect -4707 438 -4695 472
rect -4627 438 -4615 472
rect -4707 432 -4615 438
rect -4549 472 -4457 478
rect -4549 438 -4537 472
rect -4469 438 -4457 472
rect -4549 432 -4457 438
rect -4391 472 -4299 478
rect -4391 438 -4379 472
rect -4311 438 -4299 472
rect -4391 432 -4299 438
rect -4233 472 -4141 478
rect -4233 438 -4221 472
rect -4153 438 -4141 472
rect -4233 432 -4141 438
rect -4075 472 -3983 478
rect -4075 438 -4063 472
rect -3995 438 -3983 472
rect -4075 432 -3983 438
rect -3917 472 -3825 478
rect -3917 438 -3905 472
rect -3837 438 -3825 472
rect -3917 432 -3825 438
rect -3759 472 -3667 478
rect -3759 438 -3747 472
rect -3679 438 -3667 472
rect -3759 432 -3667 438
rect -3601 472 -3509 478
rect -3601 438 -3589 472
rect -3521 438 -3509 472
rect -3601 432 -3509 438
rect -3443 472 -3351 478
rect -3443 438 -3431 472
rect -3363 438 -3351 472
rect -3443 432 -3351 438
rect -3285 472 -3193 478
rect -3285 438 -3273 472
rect -3205 438 -3193 472
rect -3285 432 -3193 438
rect -3127 472 -3035 478
rect -3127 438 -3115 472
rect -3047 438 -3035 472
rect -3127 432 -3035 438
rect -2969 472 -2877 478
rect -2969 438 -2957 472
rect -2889 438 -2877 472
rect -2969 432 -2877 438
rect -2811 472 -2719 478
rect -2811 438 -2799 472
rect -2731 438 -2719 472
rect -2811 432 -2719 438
rect -2653 472 -2561 478
rect -2653 438 -2641 472
rect -2573 438 -2561 472
rect -2653 432 -2561 438
rect -2495 472 -2403 478
rect -2495 438 -2483 472
rect -2415 438 -2403 472
rect -2495 432 -2403 438
rect -2337 472 -2245 478
rect -2337 438 -2325 472
rect -2257 438 -2245 472
rect -2337 432 -2245 438
rect -2179 472 -2087 478
rect -2179 438 -2167 472
rect -2099 438 -2087 472
rect -2179 432 -2087 438
rect -2021 472 -1929 478
rect -2021 438 -2009 472
rect -1941 438 -1929 472
rect -2021 432 -1929 438
rect -1863 472 -1771 478
rect -1863 438 -1851 472
rect -1783 438 -1771 472
rect -1863 432 -1771 438
rect -1705 472 -1613 478
rect -1705 438 -1693 472
rect -1625 438 -1613 472
rect -1705 432 -1613 438
rect -1547 472 -1455 478
rect -1547 438 -1535 472
rect -1467 438 -1455 472
rect -1547 432 -1455 438
rect -1389 472 -1297 478
rect -1389 438 -1377 472
rect -1309 438 -1297 472
rect -1389 432 -1297 438
rect -1231 472 -1139 478
rect -1231 438 -1219 472
rect -1151 438 -1139 472
rect -1231 432 -1139 438
rect -1073 472 -981 478
rect -1073 438 -1061 472
rect -993 438 -981 472
rect -1073 432 -981 438
rect -915 472 -823 478
rect -915 438 -903 472
rect -835 438 -823 472
rect -915 432 -823 438
rect -757 472 -665 478
rect -757 438 -745 472
rect -677 438 -665 472
rect -757 432 -665 438
rect -599 472 -507 478
rect -599 438 -587 472
rect -519 438 -507 472
rect -599 432 -507 438
rect -441 472 -349 478
rect -441 438 -429 472
rect -361 438 -349 472
rect -441 432 -349 438
rect -283 472 -191 478
rect -283 438 -271 472
rect -203 438 -191 472
rect -283 432 -191 438
rect -125 472 -33 478
rect -125 438 -113 472
rect -45 438 -33 472
rect -125 432 -33 438
rect 33 472 125 478
rect 33 438 45 472
rect 113 438 125 472
rect 33 432 125 438
rect 191 472 283 478
rect 191 438 203 472
rect 271 438 283 472
rect 191 432 283 438
rect 349 472 441 478
rect 349 438 361 472
rect 429 438 441 472
rect 349 432 441 438
rect 507 472 599 478
rect 507 438 519 472
rect 587 438 599 472
rect 507 432 599 438
rect 665 472 757 478
rect 665 438 677 472
rect 745 438 757 472
rect 665 432 757 438
rect 823 472 915 478
rect 823 438 835 472
rect 903 438 915 472
rect 823 432 915 438
rect 981 472 1073 478
rect 981 438 993 472
rect 1061 438 1073 472
rect 981 432 1073 438
rect 1139 472 1231 478
rect 1139 438 1151 472
rect 1219 438 1231 472
rect 1139 432 1231 438
rect 1297 472 1389 478
rect 1297 438 1309 472
rect 1377 438 1389 472
rect 1297 432 1389 438
rect 1455 472 1547 478
rect 1455 438 1467 472
rect 1535 438 1547 472
rect 1455 432 1547 438
rect 1613 472 1705 478
rect 1613 438 1625 472
rect 1693 438 1705 472
rect 1613 432 1705 438
rect 1771 472 1863 478
rect 1771 438 1783 472
rect 1851 438 1863 472
rect 1771 432 1863 438
rect 1929 472 2021 478
rect 1929 438 1941 472
rect 2009 438 2021 472
rect 1929 432 2021 438
rect 2087 472 2179 478
rect 2087 438 2099 472
rect 2167 438 2179 472
rect 2087 432 2179 438
rect 2245 472 2337 478
rect 2245 438 2257 472
rect 2325 438 2337 472
rect 2245 432 2337 438
rect 2403 472 2495 478
rect 2403 438 2415 472
rect 2483 438 2495 472
rect 2403 432 2495 438
rect 2561 472 2653 478
rect 2561 438 2573 472
rect 2641 438 2653 472
rect 2561 432 2653 438
rect 2719 472 2811 478
rect 2719 438 2731 472
rect 2799 438 2811 472
rect 2719 432 2811 438
rect 2877 472 2969 478
rect 2877 438 2889 472
rect 2957 438 2969 472
rect 2877 432 2969 438
rect 3035 472 3127 478
rect 3035 438 3047 472
rect 3115 438 3127 472
rect 3035 432 3127 438
rect 3193 472 3285 478
rect 3193 438 3205 472
rect 3273 438 3285 472
rect 3193 432 3285 438
rect 3351 472 3443 478
rect 3351 438 3363 472
rect 3431 438 3443 472
rect 3351 432 3443 438
rect 3509 472 3601 478
rect 3509 438 3521 472
rect 3589 438 3601 472
rect 3509 432 3601 438
rect 3667 472 3759 478
rect 3667 438 3679 472
rect 3747 438 3759 472
rect 3667 432 3759 438
rect 3825 472 3917 478
rect 3825 438 3837 472
rect 3905 438 3917 472
rect 3825 432 3917 438
rect 3983 472 4075 478
rect 3983 438 3995 472
rect 4063 438 4075 472
rect 3983 432 4075 438
rect 4141 472 4233 478
rect 4141 438 4153 472
rect 4221 438 4233 472
rect 4141 432 4233 438
rect 4299 472 4391 478
rect 4299 438 4311 472
rect 4379 438 4391 472
rect 4299 432 4391 438
rect 4457 472 4549 478
rect 4457 438 4469 472
rect 4537 438 4549 472
rect 4457 432 4549 438
rect 4615 472 4707 478
rect 4615 438 4627 472
rect 4695 438 4707 472
rect 4615 432 4707 438
rect 4773 472 4865 478
rect 4773 438 4785 472
rect 4853 438 4865 472
rect 4773 432 4865 438
rect 4931 472 5023 478
rect 4931 438 4943 472
rect 5011 438 5023 472
rect 4931 432 5023 438
rect 5089 472 5181 478
rect 5089 438 5101 472
rect 5169 438 5181 472
rect 5089 432 5181 438
rect 5247 472 5339 478
rect 5247 438 5259 472
rect 5327 438 5339 472
rect 5247 432 5339 438
rect 5405 472 5497 478
rect 5405 438 5417 472
rect 5485 438 5497 472
rect 5405 432 5497 438
rect 5563 472 5655 478
rect 5563 438 5575 472
rect 5643 438 5655 472
rect 5563 432 5655 438
rect 5721 472 5813 478
rect 5721 438 5733 472
rect 5801 438 5813 472
rect 5721 432 5813 438
rect 5879 472 5971 478
rect 5879 438 5891 472
rect 5959 438 5971 472
rect 5879 432 5971 438
rect 6037 472 6129 478
rect 6037 438 6049 472
rect 6117 438 6129 472
rect 6037 432 6129 438
rect 6195 472 6287 478
rect 6195 438 6207 472
rect 6275 438 6287 472
rect 6195 432 6287 438
rect -6343 388 -6297 400
rect -6343 -388 -6337 388
rect -6303 -388 -6297 388
rect -6343 -400 -6297 -388
rect -6185 388 -6139 400
rect -6185 -388 -6179 388
rect -6145 -388 -6139 388
rect -6185 -400 -6139 -388
rect -6027 388 -5981 400
rect -6027 -388 -6021 388
rect -5987 -388 -5981 388
rect -6027 -400 -5981 -388
rect -5869 388 -5823 400
rect -5869 -388 -5863 388
rect -5829 -388 -5823 388
rect -5869 -400 -5823 -388
rect -5711 388 -5665 400
rect -5711 -388 -5705 388
rect -5671 -388 -5665 388
rect -5711 -400 -5665 -388
rect -5553 388 -5507 400
rect -5553 -388 -5547 388
rect -5513 -388 -5507 388
rect -5553 -400 -5507 -388
rect -5395 388 -5349 400
rect -5395 -388 -5389 388
rect -5355 -388 -5349 388
rect -5395 -400 -5349 -388
rect -5237 388 -5191 400
rect -5237 -388 -5231 388
rect -5197 -388 -5191 388
rect -5237 -400 -5191 -388
rect -5079 388 -5033 400
rect -5079 -388 -5073 388
rect -5039 -388 -5033 388
rect -5079 -400 -5033 -388
rect -4921 388 -4875 400
rect -4921 -388 -4915 388
rect -4881 -388 -4875 388
rect -4921 -400 -4875 -388
rect -4763 388 -4717 400
rect -4763 -388 -4757 388
rect -4723 -388 -4717 388
rect -4763 -400 -4717 -388
rect -4605 388 -4559 400
rect -4605 -388 -4599 388
rect -4565 -388 -4559 388
rect -4605 -400 -4559 -388
rect -4447 388 -4401 400
rect -4447 -388 -4441 388
rect -4407 -388 -4401 388
rect -4447 -400 -4401 -388
rect -4289 388 -4243 400
rect -4289 -388 -4283 388
rect -4249 -388 -4243 388
rect -4289 -400 -4243 -388
rect -4131 388 -4085 400
rect -4131 -388 -4125 388
rect -4091 -388 -4085 388
rect -4131 -400 -4085 -388
rect -3973 388 -3927 400
rect -3973 -388 -3967 388
rect -3933 -388 -3927 388
rect -3973 -400 -3927 -388
rect -3815 388 -3769 400
rect -3815 -388 -3809 388
rect -3775 -388 -3769 388
rect -3815 -400 -3769 -388
rect -3657 388 -3611 400
rect -3657 -388 -3651 388
rect -3617 -388 -3611 388
rect -3657 -400 -3611 -388
rect -3499 388 -3453 400
rect -3499 -388 -3493 388
rect -3459 -388 -3453 388
rect -3499 -400 -3453 -388
rect -3341 388 -3295 400
rect -3341 -388 -3335 388
rect -3301 -388 -3295 388
rect -3341 -400 -3295 -388
rect -3183 388 -3137 400
rect -3183 -388 -3177 388
rect -3143 -388 -3137 388
rect -3183 -400 -3137 -388
rect -3025 388 -2979 400
rect -3025 -388 -3019 388
rect -2985 -388 -2979 388
rect -3025 -400 -2979 -388
rect -2867 388 -2821 400
rect -2867 -388 -2861 388
rect -2827 -388 -2821 388
rect -2867 -400 -2821 -388
rect -2709 388 -2663 400
rect -2709 -388 -2703 388
rect -2669 -388 -2663 388
rect -2709 -400 -2663 -388
rect -2551 388 -2505 400
rect -2551 -388 -2545 388
rect -2511 -388 -2505 388
rect -2551 -400 -2505 -388
rect -2393 388 -2347 400
rect -2393 -388 -2387 388
rect -2353 -388 -2347 388
rect -2393 -400 -2347 -388
rect -2235 388 -2189 400
rect -2235 -388 -2229 388
rect -2195 -388 -2189 388
rect -2235 -400 -2189 -388
rect -2077 388 -2031 400
rect -2077 -388 -2071 388
rect -2037 -388 -2031 388
rect -2077 -400 -2031 -388
rect -1919 388 -1873 400
rect -1919 -388 -1913 388
rect -1879 -388 -1873 388
rect -1919 -400 -1873 -388
rect -1761 388 -1715 400
rect -1761 -388 -1755 388
rect -1721 -388 -1715 388
rect -1761 -400 -1715 -388
rect -1603 388 -1557 400
rect -1603 -388 -1597 388
rect -1563 -388 -1557 388
rect -1603 -400 -1557 -388
rect -1445 388 -1399 400
rect -1445 -388 -1439 388
rect -1405 -388 -1399 388
rect -1445 -400 -1399 -388
rect -1287 388 -1241 400
rect -1287 -388 -1281 388
rect -1247 -388 -1241 388
rect -1287 -400 -1241 -388
rect -1129 388 -1083 400
rect -1129 -388 -1123 388
rect -1089 -388 -1083 388
rect -1129 -400 -1083 -388
rect -971 388 -925 400
rect -971 -388 -965 388
rect -931 -388 -925 388
rect -971 -400 -925 -388
rect -813 388 -767 400
rect -813 -388 -807 388
rect -773 -388 -767 388
rect -813 -400 -767 -388
rect -655 388 -609 400
rect -655 -388 -649 388
rect -615 -388 -609 388
rect -655 -400 -609 -388
rect -497 388 -451 400
rect -497 -388 -491 388
rect -457 -388 -451 388
rect -497 -400 -451 -388
rect -339 388 -293 400
rect -339 -388 -333 388
rect -299 -388 -293 388
rect -339 -400 -293 -388
rect -181 388 -135 400
rect -181 -388 -175 388
rect -141 -388 -135 388
rect -181 -400 -135 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 135 388 181 400
rect 135 -388 141 388
rect 175 -388 181 388
rect 135 -400 181 -388
rect 293 388 339 400
rect 293 -388 299 388
rect 333 -388 339 388
rect 293 -400 339 -388
rect 451 388 497 400
rect 451 -388 457 388
rect 491 -388 497 388
rect 451 -400 497 -388
rect 609 388 655 400
rect 609 -388 615 388
rect 649 -388 655 388
rect 609 -400 655 -388
rect 767 388 813 400
rect 767 -388 773 388
rect 807 -388 813 388
rect 767 -400 813 -388
rect 925 388 971 400
rect 925 -388 931 388
rect 965 -388 971 388
rect 925 -400 971 -388
rect 1083 388 1129 400
rect 1083 -388 1089 388
rect 1123 -388 1129 388
rect 1083 -400 1129 -388
rect 1241 388 1287 400
rect 1241 -388 1247 388
rect 1281 -388 1287 388
rect 1241 -400 1287 -388
rect 1399 388 1445 400
rect 1399 -388 1405 388
rect 1439 -388 1445 388
rect 1399 -400 1445 -388
rect 1557 388 1603 400
rect 1557 -388 1563 388
rect 1597 -388 1603 388
rect 1557 -400 1603 -388
rect 1715 388 1761 400
rect 1715 -388 1721 388
rect 1755 -388 1761 388
rect 1715 -400 1761 -388
rect 1873 388 1919 400
rect 1873 -388 1879 388
rect 1913 -388 1919 388
rect 1873 -400 1919 -388
rect 2031 388 2077 400
rect 2031 -388 2037 388
rect 2071 -388 2077 388
rect 2031 -400 2077 -388
rect 2189 388 2235 400
rect 2189 -388 2195 388
rect 2229 -388 2235 388
rect 2189 -400 2235 -388
rect 2347 388 2393 400
rect 2347 -388 2353 388
rect 2387 -388 2393 388
rect 2347 -400 2393 -388
rect 2505 388 2551 400
rect 2505 -388 2511 388
rect 2545 -388 2551 388
rect 2505 -400 2551 -388
rect 2663 388 2709 400
rect 2663 -388 2669 388
rect 2703 -388 2709 388
rect 2663 -400 2709 -388
rect 2821 388 2867 400
rect 2821 -388 2827 388
rect 2861 -388 2867 388
rect 2821 -400 2867 -388
rect 2979 388 3025 400
rect 2979 -388 2985 388
rect 3019 -388 3025 388
rect 2979 -400 3025 -388
rect 3137 388 3183 400
rect 3137 -388 3143 388
rect 3177 -388 3183 388
rect 3137 -400 3183 -388
rect 3295 388 3341 400
rect 3295 -388 3301 388
rect 3335 -388 3341 388
rect 3295 -400 3341 -388
rect 3453 388 3499 400
rect 3453 -388 3459 388
rect 3493 -388 3499 388
rect 3453 -400 3499 -388
rect 3611 388 3657 400
rect 3611 -388 3617 388
rect 3651 -388 3657 388
rect 3611 -400 3657 -388
rect 3769 388 3815 400
rect 3769 -388 3775 388
rect 3809 -388 3815 388
rect 3769 -400 3815 -388
rect 3927 388 3973 400
rect 3927 -388 3933 388
rect 3967 -388 3973 388
rect 3927 -400 3973 -388
rect 4085 388 4131 400
rect 4085 -388 4091 388
rect 4125 -388 4131 388
rect 4085 -400 4131 -388
rect 4243 388 4289 400
rect 4243 -388 4249 388
rect 4283 -388 4289 388
rect 4243 -400 4289 -388
rect 4401 388 4447 400
rect 4401 -388 4407 388
rect 4441 -388 4447 388
rect 4401 -400 4447 -388
rect 4559 388 4605 400
rect 4559 -388 4565 388
rect 4599 -388 4605 388
rect 4559 -400 4605 -388
rect 4717 388 4763 400
rect 4717 -388 4723 388
rect 4757 -388 4763 388
rect 4717 -400 4763 -388
rect 4875 388 4921 400
rect 4875 -388 4881 388
rect 4915 -388 4921 388
rect 4875 -400 4921 -388
rect 5033 388 5079 400
rect 5033 -388 5039 388
rect 5073 -388 5079 388
rect 5033 -400 5079 -388
rect 5191 388 5237 400
rect 5191 -388 5197 388
rect 5231 -388 5237 388
rect 5191 -400 5237 -388
rect 5349 388 5395 400
rect 5349 -388 5355 388
rect 5389 -388 5395 388
rect 5349 -400 5395 -388
rect 5507 388 5553 400
rect 5507 -388 5513 388
rect 5547 -388 5553 388
rect 5507 -400 5553 -388
rect 5665 388 5711 400
rect 5665 -388 5671 388
rect 5705 -388 5711 388
rect 5665 -400 5711 -388
rect 5823 388 5869 400
rect 5823 -388 5829 388
rect 5863 -388 5869 388
rect 5823 -400 5869 -388
rect 5981 388 6027 400
rect 5981 -388 5987 388
rect 6021 -388 6027 388
rect 5981 -400 6027 -388
rect 6139 388 6185 400
rect 6139 -388 6145 388
rect 6179 -388 6185 388
rect 6139 -400 6185 -388
rect 6297 388 6343 400
rect 6297 -388 6303 388
rect 6337 -388 6343 388
rect 6297 -400 6343 -388
rect -6287 -438 -6195 -432
rect -6287 -472 -6275 -438
rect -6207 -472 -6195 -438
rect -6287 -478 -6195 -472
rect -6129 -438 -6037 -432
rect -6129 -472 -6117 -438
rect -6049 -472 -6037 -438
rect -6129 -478 -6037 -472
rect -5971 -438 -5879 -432
rect -5971 -472 -5959 -438
rect -5891 -472 -5879 -438
rect -5971 -478 -5879 -472
rect -5813 -438 -5721 -432
rect -5813 -472 -5801 -438
rect -5733 -472 -5721 -438
rect -5813 -478 -5721 -472
rect -5655 -438 -5563 -432
rect -5655 -472 -5643 -438
rect -5575 -472 -5563 -438
rect -5655 -478 -5563 -472
rect -5497 -438 -5405 -432
rect -5497 -472 -5485 -438
rect -5417 -472 -5405 -438
rect -5497 -478 -5405 -472
rect -5339 -438 -5247 -432
rect -5339 -472 -5327 -438
rect -5259 -472 -5247 -438
rect -5339 -478 -5247 -472
rect -5181 -438 -5089 -432
rect -5181 -472 -5169 -438
rect -5101 -472 -5089 -438
rect -5181 -478 -5089 -472
rect -5023 -438 -4931 -432
rect -5023 -472 -5011 -438
rect -4943 -472 -4931 -438
rect -5023 -478 -4931 -472
rect -4865 -438 -4773 -432
rect -4865 -472 -4853 -438
rect -4785 -472 -4773 -438
rect -4865 -478 -4773 -472
rect -4707 -438 -4615 -432
rect -4707 -472 -4695 -438
rect -4627 -472 -4615 -438
rect -4707 -478 -4615 -472
rect -4549 -438 -4457 -432
rect -4549 -472 -4537 -438
rect -4469 -472 -4457 -438
rect -4549 -478 -4457 -472
rect -4391 -438 -4299 -432
rect -4391 -472 -4379 -438
rect -4311 -472 -4299 -438
rect -4391 -478 -4299 -472
rect -4233 -438 -4141 -432
rect -4233 -472 -4221 -438
rect -4153 -472 -4141 -438
rect -4233 -478 -4141 -472
rect -4075 -438 -3983 -432
rect -4075 -472 -4063 -438
rect -3995 -472 -3983 -438
rect -4075 -478 -3983 -472
rect -3917 -438 -3825 -432
rect -3917 -472 -3905 -438
rect -3837 -472 -3825 -438
rect -3917 -478 -3825 -472
rect -3759 -438 -3667 -432
rect -3759 -472 -3747 -438
rect -3679 -472 -3667 -438
rect -3759 -478 -3667 -472
rect -3601 -438 -3509 -432
rect -3601 -472 -3589 -438
rect -3521 -472 -3509 -438
rect -3601 -478 -3509 -472
rect -3443 -438 -3351 -432
rect -3443 -472 -3431 -438
rect -3363 -472 -3351 -438
rect -3443 -478 -3351 -472
rect -3285 -438 -3193 -432
rect -3285 -472 -3273 -438
rect -3205 -472 -3193 -438
rect -3285 -478 -3193 -472
rect -3127 -438 -3035 -432
rect -3127 -472 -3115 -438
rect -3047 -472 -3035 -438
rect -3127 -478 -3035 -472
rect -2969 -438 -2877 -432
rect -2969 -472 -2957 -438
rect -2889 -472 -2877 -438
rect -2969 -478 -2877 -472
rect -2811 -438 -2719 -432
rect -2811 -472 -2799 -438
rect -2731 -472 -2719 -438
rect -2811 -478 -2719 -472
rect -2653 -438 -2561 -432
rect -2653 -472 -2641 -438
rect -2573 -472 -2561 -438
rect -2653 -478 -2561 -472
rect -2495 -438 -2403 -432
rect -2495 -472 -2483 -438
rect -2415 -472 -2403 -438
rect -2495 -478 -2403 -472
rect -2337 -438 -2245 -432
rect -2337 -472 -2325 -438
rect -2257 -472 -2245 -438
rect -2337 -478 -2245 -472
rect -2179 -438 -2087 -432
rect -2179 -472 -2167 -438
rect -2099 -472 -2087 -438
rect -2179 -478 -2087 -472
rect -2021 -438 -1929 -432
rect -2021 -472 -2009 -438
rect -1941 -472 -1929 -438
rect -2021 -478 -1929 -472
rect -1863 -438 -1771 -432
rect -1863 -472 -1851 -438
rect -1783 -472 -1771 -438
rect -1863 -478 -1771 -472
rect -1705 -438 -1613 -432
rect -1705 -472 -1693 -438
rect -1625 -472 -1613 -438
rect -1705 -478 -1613 -472
rect -1547 -438 -1455 -432
rect -1547 -472 -1535 -438
rect -1467 -472 -1455 -438
rect -1547 -478 -1455 -472
rect -1389 -438 -1297 -432
rect -1389 -472 -1377 -438
rect -1309 -472 -1297 -438
rect -1389 -478 -1297 -472
rect -1231 -438 -1139 -432
rect -1231 -472 -1219 -438
rect -1151 -472 -1139 -438
rect -1231 -478 -1139 -472
rect -1073 -438 -981 -432
rect -1073 -472 -1061 -438
rect -993 -472 -981 -438
rect -1073 -478 -981 -472
rect -915 -438 -823 -432
rect -915 -472 -903 -438
rect -835 -472 -823 -438
rect -915 -478 -823 -472
rect -757 -438 -665 -432
rect -757 -472 -745 -438
rect -677 -472 -665 -438
rect -757 -478 -665 -472
rect -599 -438 -507 -432
rect -599 -472 -587 -438
rect -519 -472 -507 -438
rect -599 -478 -507 -472
rect -441 -438 -349 -432
rect -441 -472 -429 -438
rect -361 -472 -349 -438
rect -441 -478 -349 -472
rect -283 -438 -191 -432
rect -283 -472 -271 -438
rect -203 -472 -191 -438
rect -283 -478 -191 -472
rect -125 -438 -33 -432
rect -125 -472 -113 -438
rect -45 -472 -33 -438
rect -125 -478 -33 -472
rect 33 -438 125 -432
rect 33 -472 45 -438
rect 113 -472 125 -438
rect 33 -478 125 -472
rect 191 -438 283 -432
rect 191 -472 203 -438
rect 271 -472 283 -438
rect 191 -478 283 -472
rect 349 -438 441 -432
rect 349 -472 361 -438
rect 429 -472 441 -438
rect 349 -478 441 -472
rect 507 -438 599 -432
rect 507 -472 519 -438
rect 587 -472 599 -438
rect 507 -478 599 -472
rect 665 -438 757 -432
rect 665 -472 677 -438
rect 745 -472 757 -438
rect 665 -478 757 -472
rect 823 -438 915 -432
rect 823 -472 835 -438
rect 903 -472 915 -438
rect 823 -478 915 -472
rect 981 -438 1073 -432
rect 981 -472 993 -438
rect 1061 -472 1073 -438
rect 981 -478 1073 -472
rect 1139 -438 1231 -432
rect 1139 -472 1151 -438
rect 1219 -472 1231 -438
rect 1139 -478 1231 -472
rect 1297 -438 1389 -432
rect 1297 -472 1309 -438
rect 1377 -472 1389 -438
rect 1297 -478 1389 -472
rect 1455 -438 1547 -432
rect 1455 -472 1467 -438
rect 1535 -472 1547 -438
rect 1455 -478 1547 -472
rect 1613 -438 1705 -432
rect 1613 -472 1625 -438
rect 1693 -472 1705 -438
rect 1613 -478 1705 -472
rect 1771 -438 1863 -432
rect 1771 -472 1783 -438
rect 1851 -472 1863 -438
rect 1771 -478 1863 -472
rect 1929 -438 2021 -432
rect 1929 -472 1941 -438
rect 2009 -472 2021 -438
rect 1929 -478 2021 -472
rect 2087 -438 2179 -432
rect 2087 -472 2099 -438
rect 2167 -472 2179 -438
rect 2087 -478 2179 -472
rect 2245 -438 2337 -432
rect 2245 -472 2257 -438
rect 2325 -472 2337 -438
rect 2245 -478 2337 -472
rect 2403 -438 2495 -432
rect 2403 -472 2415 -438
rect 2483 -472 2495 -438
rect 2403 -478 2495 -472
rect 2561 -438 2653 -432
rect 2561 -472 2573 -438
rect 2641 -472 2653 -438
rect 2561 -478 2653 -472
rect 2719 -438 2811 -432
rect 2719 -472 2731 -438
rect 2799 -472 2811 -438
rect 2719 -478 2811 -472
rect 2877 -438 2969 -432
rect 2877 -472 2889 -438
rect 2957 -472 2969 -438
rect 2877 -478 2969 -472
rect 3035 -438 3127 -432
rect 3035 -472 3047 -438
rect 3115 -472 3127 -438
rect 3035 -478 3127 -472
rect 3193 -438 3285 -432
rect 3193 -472 3205 -438
rect 3273 -472 3285 -438
rect 3193 -478 3285 -472
rect 3351 -438 3443 -432
rect 3351 -472 3363 -438
rect 3431 -472 3443 -438
rect 3351 -478 3443 -472
rect 3509 -438 3601 -432
rect 3509 -472 3521 -438
rect 3589 -472 3601 -438
rect 3509 -478 3601 -472
rect 3667 -438 3759 -432
rect 3667 -472 3679 -438
rect 3747 -472 3759 -438
rect 3667 -478 3759 -472
rect 3825 -438 3917 -432
rect 3825 -472 3837 -438
rect 3905 -472 3917 -438
rect 3825 -478 3917 -472
rect 3983 -438 4075 -432
rect 3983 -472 3995 -438
rect 4063 -472 4075 -438
rect 3983 -478 4075 -472
rect 4141 -438 4233 -432
rect 4141 -472 4153 -438
rect 4221 -472 4233 -438
rect 4141 -478 4233 -472
rect 4299 -438 4391 -432
rect 4299 -472 4311 -438
rect 4379 -472 4391 -438
rect 4299 -478 4391 -472
rect 4457 -438 4549 -432
rect 4457 -472 4469 -438
rect 4537 -472 4549 -438
rect 4457 -478 4549 -472
rect 4615 -438 4707 -432
rect 4615 -472 4627 -438
rect 4695 -472 4707 -438
rect 4615 -478 4707 -472
rect 4773 -438 4865 -432
rect 4773 -472 4785 -438
rect 4853 -472 4865 -438
rect 4773 -478 4865 -472
rect 4931 -438 5023 -432
rect 4931 -472 4943 -438
rect 5011 -472 5023 -438
rect 4931 -478 5023 -472
rect 5089 -438 5181 -432
rect 5089 -472 5101 -438
rect 5169 -472 5181 -438
rect 5089 -478 5181 -472
rect 5247 -438 5339 -432
rect 5247 -472 5259 -438
rect 5327 -472 5339 -438
rect 5247 -478 5339 -472
rect 5405 -438 5497 -432
rect 5405 -472 5417 -438
rect 5485 -472 5497 -438
rect 5405 -478 5497 -472
rect 5563 -438 5655 -432
rect 5563 -472 5575 -438
rect 5643 -472 5655 -438
rect 5563 -478 5655 -472
rect 5721 -438 5813 -432
rect 5721 -472 5733 -438
rect 5801 -472 5813 -438
rect 5721 -478 5813 -472
rect 5879 -438 5971 -432
rect 5879 -472 5891 -438
rect 5959 -472 5971 -438
rect 5879 -478 5971 -472
rect 6037 -438 6129 -432
rect 6037 -472 6049 -438
rect 6117 -472 6129 -438
rect 6037 -478 6129 -472
rect 6195 -438 6287 -432
rect 6195 -472 6207 -438
rect 6275 -472 6287 -438
rect 6195 -478 6287 -472
rect -6343 -522 -6297 -510
rect -6343 -1298 -6337 -522
rect -6303 -1298 -6297 -522
rect -6343 -1310 -6297 -1298
rect -6185 -522 -6139 -510
rect -6185 -1298 -6179 -522
rect -6145 -1298 -6139 -522
rect -6185 -1310 -6139 -1298
rect -6027 -522 -5981 -510
rect -6027 -1298 -6021 -522
rect -5987 -1298 -5981 -522
rect -6027 -1310 -5981 -1298
rect -5869 -522 -5823 -510
rect -5869 -1298 -5863 -522
rect -5829 -1298 -5823 -522
rect -5869 -1310 -5823 -1298
rect -5711 -522 -5665 -510
rect -5711 -1298 -5705 -522
rect -5671 -1298 -5665 -522
rect -5711 -1310 -5665 -1298
rect -5553 -522 -5507 -510
rect -5553 -1298 -5547 -522
rect -5513 -1298 -5507 -522
rect -5553 -1310 -5507 -1298
rect -5395 -522 -5349 -510
rect -5395 -1298 -5389 -522
rect -5355 -1298 -5349 -522
rect -5395 -1310 -5349 -1298
rect -5237 -522 -5191 -510
rect -5237 -1298 -5231 -522
rect -5197 -1298 -5191 -522
rect -5237 -1310 -5191 -1298
rect -5079 -522 -5033 -510
rect -5079 -1298 -5073 -522
rect -5039 -1298 -5033 -522
rect -5079 -1310 -5033 -1298
rect -4921 -522 -4875 -510
rect -4921 -1298 -4915 -522
rect -4881 -1298 -4875 -522
rect -4921 -1310 -4875 -1298
rect -4763 -522 -4717 -510
rect -4763 -1298 -4757 -522
rect -4723 -1298 -4717 -522
rect -4763 -1310 -4717 -1298
rect -4605 -522 -4559 -510
rect -4605 -1298 -4599 -522
rect -4565 -1298 -4559 -522
rect -4605 -1310 -4559 -1298
rect -4447 -522 -4401 -510
rect -4447 -1298 -4441 -522
rect -4407 -1298 -4401 -522
rect -4447 -1310 -4401 -1298
rect -4289 -522 -4243 -510
rect -4289 -1298 -4283 -522
rect -4249 -1298 -4243 -522
rect -4289 -1310 -4243 -1298
rect -4131 -522 -4085 -510
rect -4131 -1298 -4125 -522
rect -4091 -1298 -4085 -522
rect -4131 -1310 -4085 -1298
rect -3973 -522 -3927 -510
rect -3973 -1298 -3967 -522
rect -3933 -1298 -3927 -522
rect -3973 -1310 -3927 -1298
rect -3815 -522 -3769 -510
rect -3815 -1298 -3809 -522
rect -3775 -1298 -3769 -522
rect -3815 -1310 -3769 -1298
rect -3657 -522 -3611 -510
rect -3657 -1298 -3651 -522
rect -3617 -1298 -3611 -522
rect -3657 -1310 -3611 -1298
rect -3499 -522 -3453 -510
rect -3499 -1298 -3493 -522
rect -3459 -1298 -3453 -522
rect -3499 -1310 -3453 -1298
rect -3341 -522 -3295 -510
rect -3341 -1298 -3335 -522
rect -3301 -1298 -3295 -522
rect -3341 -1310 -3295 -1298
rect -3183 -522 -3137 -510
rect -3183 -1298 -3177 -522
rect -3143 -1298 -3137 -522
rect -3183 -1310 -3137 -1298
rect -3025 -522 -2979 -510
rect -3025 -1298 -3019 -522
rect -2985 -1298 -2979 -522
rect -3025 -1310 -2979 -1298
rect -2867 -522 -2821 -510
rect -2867 -1298 -2861 -522
rect -2827 -1298 -2821 -522
rect -2867 -1310 -2821 -1298
rect -2709 -522 -2663 -510
rect -2709 -1298 -2703 -522
rect -2669 -1298 -2663 -522
rect -2709 -1310 -2663 -1298
rect -2551 -522 -2505 -510
rect -2551 -1298 -2545 -522
rect -2511 -1298 -2505 -522
rect -2551 -1310 -2505 -1298
rect -2393 -522 -2347 -510
rect -2393 -1298 -2387 -522
rect -2353 -1298 -2347 -522
rect -2393 -1310 -2347 -1298
rect -2235 -522 -2189 -510
rect -2235 -1298 -2229 -522
rect -2195 -1298 -2189 -522
rect -2235 -1310 -2189 -1298
rect -2077 -522 -2031 -510
rect -2077 -1298 -2071 -522
rect -2037 -1298 -2031 -522
rect -2077 -1310 -2031 -1298
rect -1919 -522 -1873 -510
rect -1919 -1298 -1913 -522
rect -1879 -1298 -1873 -522
rect -1919 -1310 -1873 -1298
rect -1761 -522 -1715 -510
rect -1761 -1298 -1755 -522
rect -1721 -1298 -1715 -522
rect -1761 -1310 -1715 -1298
rect -1603 -522 -1557 -510
rect -1603 -1298 -1597 -522
rect -1563 -1298 -1557 -522
rect -1603 -1310 -1557 -1298
rect -1445 -522 -1399 -510
rect -1445 -1298 -1439 -522
rect -1405 -1298 -1399 -522
rect -1445 -1310 -1399 -1298
rect -1287 -522 -1241 -510
rect -1287 -1298 -1281 -522
rect -1247 -1298 -1241 -522
rect -1287 -1310 -1241 -1298
rect -1129 -522 -1083 -510
rect -1129 -1298 -1123 -522
rect -1089 -1298 -1083 -522
rect -1129 -1310 -1083 -1298
rect -971 -522 -925 -510
rect -971 -1298 -965 -522
rect -931 -1298 -925 -522
rect -971 -1310 -925 -1298
rect -813 -522 -767 -510
rect -813 -1298 -807 -522
rect -773 -1298 -767 -522
rect -813 -1310 -767 -1298
rect -655 -522 -609 -510
rect -655 -1298 -649 -522
rect -615 -1298 -609 -522
rect -655 -1310 -609 -1298
rect -497 -522 -451 -510
rect -497 -1298 -491 -522
rect -457 -1298 -451 -522
rect -497 -1310 -451 -1298
rect -339 -522 -293 -510
rect -339 -1298 -333 -522
rect -299 -1298 -293 -522
rect -339 -1310 -293 -1298
rect -181 -522 -135 -510
rect -181 -1298 -175 -522
rect -141 -1298 -135 -522
rect -181 -1310 -135 -1298
rect -23 -522 23 -510
rect -23 -1298 -17 -522
rect 17 -1298 23 -522
rect -23 -1310 23 -1298
rect 135 -522 181 -510
rect 135 -1298 141 -522
rect 175 -1298 181 -522
rect 135 -1310 181 -1298
rect 293 -522 339 -510
rect 293 -1298 299 -522
rect 333 -1298 339 -522
rect 293 -1310 339 -1298
rect 451 -522 497 -510
rect 451 -1298 457 -522
rect 491 -1298 497 -522
rect 451 -1310 497 -1298
rect 609 -522 655 -510
rect 609 -1298 615 -522
rect 649 -1298 655 -522
rect 609 -1310 655 -1298
rect 767 -522 813 -510
rect 767 -1298 773 -522
rect 807 -1298 813 -522
rect 767 -1310 813 -1298
rect 925 -522 971 -510
rect 925 -1298 931 -522
rect 965 -1298 971 -522
rect 925 -1310 971 -1298
rect 1083 -522 1129 -510
rect 1083 -1298 1089 -522
rect 1123 -1298 1129 -522
rect 1083 -1310 1129 -1298
rect 1241 -522 1287 -510
rect 1241 -1298 1247 -522
rect 1281 -1298 1287 -522
rect 1241 -1310 1287 -1298
rect 1399 -522 1445 -510
rect 1399 -1298 1405 -522
rect 1439 -1298 1445 -522
rect 1399 -1310 1445 -1298
rect 1557 -522 1603 -510
rect 1557 -1298 1563 -522
rect 1597 -1298 1603 -522
rect 1557 -1310 1603 -1298
rect 1715 -522 1761 -510
rect 1715 -1298 1721 -522
rect 1755 -1298 1761 -522
rect 1715 -1310 1761 -1298
rect 1873 -522 1919 -510
rect 1873 -1298 1879 -522
rect 1913 -1298 1919 -522
rect 1873 -1310 1919 -1298
rect 2031 -522 2077 -510
rect 2031 -1298 2037 -522
rect 2071 -1298 2077 -522
rect 2031 -1310 2077 -1298
rect 2189 -522 2235 -510
rect 2189 -1298 2195 -522
rect 2229 -1298 2235 -522
rect 2189 -1310 2235 -1298
rect 2347 -522 2393 -510
rect 2347 -1298 2353 -522
rect 2387 -1298 2393 -522
rect 2347 -1310 2393 -1298
rect 2505 -522 2551 -510
rect 2505 -1298 2511 -522
rect 2545 -1298 2551 -522
rect 2505 -1310 2551 -1298
rect 2663 -522 2709 -510
rect 2663 -1298 2669 -522
rect 2703 -1298 2709 -522
rect 2663 -1310 2709 -1298
rect 2821 -522 2867 -510
rect 2821 -1298 2827 -522
rect 2861 -1298 2867 -522
rect 2821 -1310 2867 -1298
rect 2979 -522 3025 -510
rect 2979 -1298 2985 -522
rect 3019 -1298 3025 -522
rect 2979 -1310 3025 -1298
rect 3137 -522 3183 -510
rect 3137 -1298 3143 -522
rect 3177 -1298 3183 -522
rect 3137 -1310 3183 -1298
rect 3295 -522 3341 -510
rect 3295 -1298 3301 -522
rect 3335 -1298 3341 -522
rect 3295 -1310 3341 -1298
rect 3453 -522 3499 -510
rect 3453 -1298 3459 -522
rect 3493 -1298 3499 -522
rect 3453 -1310 3499 -1298
rect 3611 -522 3657 -510
rect 3611 -1298 3617 -522
rect 3651 -1298 3657 -522
rect 3611 -1310 3657 -1298
rect 3769 -522 3815 -510
rect 3769 -1298 3775 -522
rect 3809 -1298 3815 -522
rect 3769 -1310 3815 -1298
rect 3927 -522 3973 -510
rect 3927 -1298 3933 -522
rect 3967 -1298 3973 -522
rect 3927 -1310 3973 -1298
rect 4085 -522 4131 -510
rect 4085 -1298 4091 -522
rect 4125 -1298 4131 -522
rect 4085 -1310 4131 -1298
rect 4243 -522 4289 -510
rect 4243 -1298 4249 -522
rect 4283 -1298 4289 -522
rect 4243 -1310 4289 -1298
rect 4401 -522 4447 -510
rect 4401 -1298 4407 -522
rect 4441 -1298 4447 -522
rect 4401 -1310 4447 -1298
rect 4559 -522 4605 -510
rect 4559 -1298 4565 -522
rect 4599 -1298 4605 -522
rect 4559 -1310 4605 -1298
rect 4717 -522 4763 -510
rect 4717 -1298 4723 -522
rect 4757 -1298 4763 -522
rect 4717 -1310 4763 -1298
rect 4875 -522 4921 -510
rect 4875 -1298 4881 -522
rect 4915 -1298 4921 -522
rect 4875 -1310 4921 -1298
rect 5033 -522 5079 -510
rect 5033 -1298 5039 -522
rect 5073 -1298 5079 -522
rect 5033 -1310 5079 -1298
rect 5191 -522 5237 -510
rect 5191 -1298 5197 -522
rect 5231 -1298 5237 -522
rect 5191 -1310 5237 -1298
rect 5349 -522 5395 -510
rect 5349 -1298 5355 -522
rect 5389 -1298 5395 -522
rect 5349 -1310 5395 -1298
rect 5507 -522 5553 -510
rect 5507 -1298 5513 -522
rect 5547 -1298 5553 -522
rect 5507 -1310 5553 -1298
rect 5665 -522 5711 -510
rect 5665 -1298 5671 -522
rect 5705 -1298 5711 -522
rect 5665 -1310 5711 -1298
rect 5823 -522 5869 -510
rect 5823 -1298 5829 -522
rect 5863 -1298 5869 -522
rect 5823 -1310 5869 -1298
rect 5981 -522 6027 -510
rect 5981 -1298 5987 -522
rect 6021 -1298 6027 -522
rect 5981 -1310 6027 -1298
rect 6139 -522 6185 -510
rect 6139 -1298 6145 -522
rect 6179 -1298 6185 -522
rect 6139 -1310 6185 -1298
rect 6297 -522 6343 -510
rect 6297 -1298 6303 -522
rect 6337 -1298 6343 -522
rect 6297 -1310 6343 -1298
rect -6287 -1348 -6195 -1342
rect -6287 -1382 -6275 -1348
rect -6207 -1382 -6195 -1348
rect -6287 -1388 -6195 -1382
rect -6129 -1348 -6037 -1342
rect -6129 -1382 -6117 -1348
rect -6049 -1382 -6037 -1348
rect -6129 -1388 -6037 -1382
rect -5971 -1348 -5879 -1342
rect -5971 -1382 -5959 -1348
rect -5891 -1382 -5879 -1348
rect -5971 -1388 -5879 -1382
rect -5813 -1348 -5721 -1342
rect -5813 -1382 -5801 -1348
rect -5733 -1382 -5721 -1348
rect -5813 -1388 -5721 -1382
rect -5655 -1348 -5563 -1342
rect -5655 -1382 -5643 -1348
rect -5575 -1382 -5563 -1348
rect -5655 -1388 -5563 -1382
rect -5497 -1348 -5405 -1342
rect -5497 -1382 -5485 -1348
rect -5417 -1382 -5405 -1348
rect -5497 -1388 -5405 -1382
rect -5339 -1348 -5247 -1342
rect -5339 -1382 -5327 -1348
rect -5259 -1382 -5247 -1348
rect -5339 -1388 -5247 -1382
rect -5181 -1348 -5089 -1342
rect -5181 -1382 -5169 -1348
rect -5101 -1382 -5089 -1348
rect -5181 -1388 -5089 -1382
rect -5023 -1348 -4931 -1342
rect -5023 -1382 -5011 -1348
rect -4943 -1382 -4931 -1348
rect -5023 -1388 -4931 -1382
rect -4865 -1348 -4773 -1342
rect -4865 -1382 -4853 -1348
rect -4785 -1382 -4773 -1348
rect -4865 -1388 -4773 -1382
rect -4707 -1348 -4615 -1342
rect -4707 -1382 -4695 -1348
rect -4627 -1382 -4615 -1348
rect -4707 -1388 -4615 -1382
rect -4549 -1348 -4457 -1342
rect -4549 -1382 -4537 -1348
rect -4469 -1382 -4457 -1348
rect -4549 -1388 -4457 -1382
rect -4391 -1348 -4299 -1342
rect -4391 -1382 -4379 -1348
rect -4311 -1382 -4299 -1348
rect -4391 -1388 -4299 -1382
rect -4233 -1348 -4141 -1342
rect -4233 -1382 -4221 -1348
rect -4153 -1382 -4141 -1348
rect -4233 -1388 -4141 -1382
rect -4075 -1348 -3983 -1342
rect -4075 -1382 -4063 -1348
rect -3995 -1382 -3983 -1348
rect -4075 -1388 -3983 -1382
rect -3917 -1348 -3825 -1342
rect -3917 -1382 -3905 -1348
rect -3837 -1382 -3825 -1348
rect -3917 -1388 -3825 -1382
rect -3759 -1348 -3667 -1342
rect -3759 -1382 -3747 -1348
rect -3679 -1382 -3667 -1348
rect -3759 -1388 -3667 -1382
rect -3601 -1348 -3509 -1342
rect -3601 -1382 -3589 -1348
rect -3521 -1382 -3509 -1348
rect -3601 -1388 -3509 -1382
rect -3443 -1348 -3351 -1342
rect -3443 -1382 -3431 -1348
rect -3363 -1382 -3351 -1348
rect -3443 -1388 -3351 -1382
rect -3285 -1348 -3193 -1342
rect -3285 -1382 -3273 -1348
rect -3205 -1382 -3193 -1348
rect -3285 -1388 -3193 -1382
rect -3127 -1348 -3035 -1342
rect -3127 -1382 -3115 -1348
rect -3047 -1382 -3035 -1348
rect -3127 -1388 -3035 -1382
rect -2969 -1348 -2877 -1342
rect -2969 -1382 -2957 -1348
rect -2889 -1382 -2877 -1348
rect -2969 -1388 -2877 -1382
rect -2811 -1348 -2719 -1342
rect -2811 -1382 -2799 -1348
rect -2731 -1382 -2719 -1348
rect -2811 -1388 -2719 -1382
rect -2653 -1348 -2561 -1342
rect -2653 -1382 -2641 -1348
rect -2573 -1382 -2561 -1348
rect -2653 -1388 -2561 -1382
rect -2495 -1348 -2403 -1342
rect -2495 -1382 -2483 -1348
rect -2415 -1382 -2403 -1348
rect -2495 -1388 -2403 -1382
rect -2337 -1348 -2245 -1342
rect -2337 -1382 -2325 -1348
rect -2257 -1382 -2245 -1348
rect -2337 -1388 -2245 -1382
rect -2179 -1348 -2087 -1342
rect -2179 -1382 -2167 -1348
rect -2099 -1382 -2087 -1348
rect -2179 -1388 -2087 -1382
rect -2021 -1348 -1929 -1342
rect -2021 -1382 -2009 -1348
rect -1941 -1382 -1929 -1348
rect -2021 -1388 -1929 -1382
rect -1863 -1348 -1771 -1342
rect -1863 -1382 -1851 -1348
rect -1783 -1382 -1771 -1348
rect -1863 -1388 -1771 -1382
rect -1705 -1348 -1613 -1342
rect -1705 -1382 -1693 -1348
rect -1625 -1382 -1613 -1348
rect -1705 -1388 -1613 -1382
rect -1547 -1348 -1455 -1342
rect -1547 -1382 -1535 -1348
rect -1467 -1382 -1455 -1348
rect -1547 -1388 -1455 -1382
rect -1389 -1348 -1297 -1342
rect -1389 -1382 -1377 -1348
rect -1309 -1382 -1297 -1348
rect -1389 -1388 -1297 -1382
rect -1231 -1348 -1139 -1342
rect -1231 -1382 -1219 -1348
rect -1151 -1382 -1139 -1348
rect -1231 -1388 -1139 -1382
rect -1073 -1348 -981 -1342
rect -1073 -1382 -1061 -1348
rect -993 -1382 -981 -1348
rect -1073 -1388 -981 -1382
rect -915 -1348 -823 -1342
rect -915 -1382 -903 -1348
rect -835 -1382 -823 -1348
rect -915 -1388 -823 -1382
rect -757 -1348 -665 -1342
rect -757 -1382 -745 -1348
rect -677 -1382 -665 -1348
rect -757 -1388 -665 -1382
rect -599 -1348 -507 -1342
rect -599 -1382 -587 -1348
rect -519 -1382 -507 -1348
rect -599 -1388 -507 -1382
rect -441 -1348 -349 -1342
rect -441 -1382 -429 -1348
rect -361 -1382 -349 -1348
rect -441 -1388 -349 -1382
rect -283 -1348 -191 -1342
rect -283 -1382 -271 -1348
rect -203 -1382 -191 -1348
rect -283 -1388 -191 -1382
rect -125 -1348 -33 -1342
rect -125 -1382 -113 -1348
rect -45 -1382 -33 -1348
rect -125 -1388 -33 -1382
rect 33 -1348 125 -1342
rect 33 -1382 45 -1348
rect 113 -1382 125 -1348
rect 33 -1388 125 -1382
rect 191 -1348 283 -1342
rect 191 -1382 203 -1348
rect 271 -1382 283 -1348
rect 191 -1388 283 -1382
rect 349 -1348 441 -1342
rect 349 -1382 361 -1348
rect 429 -1382 441 -1348
rect 349 -1388 441 -1382
rect 507 -1348 599 -1342
rect 507 -1382 519 -1348
rect 587 -1382 599 -1348
rect 507 -1388 599 -1382
rect 665 -1348 757 -1342
rect 665 -1382 677 -1348
rect 745 -1382 757 -1348
rect 665 -1388 757 -1382
rect 823 -1348 915 -1342
rect 823 -1382 835 -1348
rect 903 -1382 915 -1348
rect 823 -1388 915 -1382
rect 981 -1348 1073 -1342
rect 981 -1382 993 -1348
rect 1061 -1382 1073 -1348
rect 981 -1388 1073 -1382
rect 1139 -1348 1231 -1342
rect 1139 -1382 1151 -1348
rect 1219 -1382 1231 -1348
rect 1139 -1388 1231 -1382
rect 1297 -1348 1389 -1342
rect 1297 -1382 1309 -1348
rect 1377 -1382 1389 -1348
rect 1297 -1388 1389 -1382
rect 1455 -1348 1547 -1342
rect 1455 -1382 1467 -1348
rect 1535 -1382 1547 -1348
rect 1455 -1388 1547 -1382
rect 1613 -1348 1705 -1342
rect 1613 -1382 1625 -1348
rect 1693 -1382 1705 -1348
rect 1613 -1388 1705 -1382
rect 1771 -1348 1863 -1342
rect 1771 -1382 1783 -1348
rect 1851 -1382 1863 -1348
rect 1771 -1388 1863 -1382
rect 1929 -1348 2021 -1342
rect 1929 -1382 1941 -1348
rect 2009 -1382 2021 -1348
rect 1929 -1388 2021 -1382
rect 2087 -1348 2179 -1342
rect 2087 -1382 2099 -1348
rect 2167 -1382 2179 -1348
rect 2087 -1388 2179 -1382
rect 2245 -1348 2337 -1342
rect 2245 -1382 2257 -1348
rect 2325 -1382 2337 -1348
rect 2245 -1388 2337 -1382
rect 2403 -1348 2495 -1342
rect 2403 -1382 2415 -1348
rect 2483 -1382 2495 -1348
rect 2403 -1388 2495 -1382
rect 2561 -1348 2653 -1342
rect 2561 -1382 2573 -1348
rect 2641 -1382 2653 -1348
rect 2561 -1388 2653 -1382
rect 2719 -1348 2811 -1342
rect 2719 -1382 2731 -1348
rect 2799 -1382 2811 -1348
rect 2719 -1388 2811 -1382
rect 2877 -1348 2969 -1342
rect 2877 -1382 2889 -1348
rect 2957 -1382 2969 -1348
rect 2877 -1388 2969 -1382
rect 3035 -1348 3127 -1342
rect 3035 -1382 3047 -1348
rect 3115 -1382 3127 -1348
rect 3035 -1388 3127 -1382
rect 3193 -1348 3285 -1342
rect 3193 -1382 3205 -1348
rect 3273 -1382 3285 -1348
rect 3193 -1388 3285 -1382
rect 3351 -1348 3443 -1342
rect 3351 -1382 3363 -1348
rect 3431 -1382 3443 -1348
rect 3351 -1388 3443 -1382
rect 3509 -1348 3601 -1342
rect 3509 -1382 3521 -1348
rect 3589 -1382 3601 -1348
rect 3509 -1388 3601 -1382
rect 3667 -1348 3759 -1342
rect 3667 -1382 3679 -1348
rect 3747 -1382 3759 -1348
rect 3667 -1388 3759 -1382
rect 3825 -1348 3917 -1342
rect 3825 -1382 3837 -1348
rect 3905 -1382 3917 -1348
rect 3825 -1388 3917 -1382
rect 3983 -1348 4075 -1342
rect 3983 -1382 3995 -1348
rect 4063 -1382 4075 -1348
rect 3983 -1388 4075 -1382
rect 4141 -1348 4233 -1342
rect 4141 -1382 4153 -1348
rect 4221 -1382 4233 -1348
rect 4141 -1388 4233 -1382
rect 4299 -1348 4391 -1342
rect 4299 -1382 4311 -1348
rect 4379 -1382 4391 -1348
rect 4299 -1388 4391 -1382
rect 4457 -1348 4549 -1342
rect 4457 -1382 4469 -1348
rect 4537 -1382 4549 -1348
rect 4457 -1388 4549 -1382
rect 4615 -1348 4707 -1342
rect 4615 -1382 4627 -1348
rect 4695 -1382 4707 -1348
rect 4615 -1388 4707 -1382
rect 4773 -1348 4865 -1342
rect 4773 -1382 4785 -1348
rect 4853 -1382 4865 -1348
rect 4773 -1388 4865 -1382
rect 4931 -1348 5023 -1342
rect 4931 -1382 4943 -1348
rect 5011 -1382 5023 -1348
rect 4931 -1388 5023 -1382
rect 5089 -1348 5181 -1342
rect 5089 -1382 5101 -1348
rect 5169 -1382 5181 -1348
rect 5089 -1388 5181 -1382
rect 5247 -1348 5339 -1342
rect 5247 -1382 5259 -1348
rect 5327 -1382 5339 -1348
rect 5247 -1388 5339 -1382
rect 5405 -1348 5497 -1342
rect 5405 -1382 5417 -1348
rect 5485 -1382 5497 -1348
rect 5405 -1388 5497 -1382
rect 5563 -1348 5655 -1342
rect 5563 -1382 5575 -1348
rect 5643 -1382 5655 -1348
rect 5563 -1388 5655 -1382
rect 5721 -1348 5813 -1342
rect 5721 -1382 5733 -1348
rect 5801 -1382 5813 -1348
rect 5721 -1388 5813 -1382
rect 5879 -1348 5971 -1342
rect 5879 -1382 5891 -1348
rect 5959 -1382 5971 -1348
rect 5879 -1388 5971 -1382
rect 6037 -1348 6129 -1342
rect 6037 -1382 6049 -1348
rect 6117 -1382 6129 -1348
rect 6037 -1388 6129 -1382
rect 6195 -1348 6287 -1342
rect 6195 -1382 6207 -1348
rect 6275 -1382 6287 -1348
rect 6195 -1388 6287 -1382
rect -6343 -1432 -6297 -1420
rect -6343 -2208 -6337 -1432
rect -6303 -2208 -6297 -1432
rect -6343 -2220 -6297 -2208
rect -6185 -1432 -6139 -1420
rect -6185 -2208 -6179 -1432
rect -6145 -2208 -6139 -1432
rect -6185 -2220 -6139 -2208
rect -6027 -1432 -5981 -1420
rect -6027 -2208 -6021 -1432
rect -5987 -2208 -5981 -1432
rect -6027 -2220 -5981 -2208
rect -5869 -1432 -5823 -1420
rect -5869 -2208 -5863 -1432
rect -5829 -2208 -5823 -1432
rect -5869 -2220 -5823 -2208
rect -5711 -1432 -5665 -1420
rect -5711 -2208 -5705 -1432
rect -5671 -2208 -5665 -1432
rect -5711 -2220 -5665 -2208
rect -5553 -1432 -5507 -1420
rect -5553 -2208 -5547 -1432
rect -5513 -2208 -5507 -1432
rect -5553 -2220 -5507 -2208
rect -5395 -1432 -5349 -1420
rect -5395 -2208 -5389 -1432
rect -5355 -2208 -5349 -1432
rect -5395 -2220 -5349 -2208
rect -5237 -1432 -5191 -1420
rect -5237 -2208 -5231 -1432
rect -5197 -2208 -5191 -1432
rect -5237 -2220 -5191 -2208
rect -5079 -1432 -5033 -1420
rect -5079 -2208 -5073 -1432
rect -5039 -2208 -5033 -1432
rect -5079 -2220 -5033 -2208
rect -4921 -1432 -4875 -1420
rect -4921 -2208 -4915 -1432
rect -4881 -2208 -4875 -1432
rect -4921 -2220 -4875 -2208
rect -4763 -1432 -4717 -1420
rect -4763 -2208 -4757 -1432
rect -4723 -2208 -4717 -1432
rect -4763 -2220 -4717 -2208
rect -4605 -1432 -4559 -1420
rect -4605 -2208 -4599 -1432
rect -4565 -2208 -4559 -1432
rect -4605 -2220 -4559 -2208
rect -4447 -1432 -4401 -1420
rect -4447 -2208 -4441 -1432
rect -4407 -2208 -4401 -1432
rect -4447 -2220 -4401 -2208
rect -4289 -1432 -4243 -1420
rect -4289 -2208 -4283 -1432
rect -4249 -2208 -4243 -1432
rect -4289 -2220 -4243 -2208
rect -4131 -1432 -4085 -1420
rect -4131 -2208 -4125 -1432
rect -4091 -2208 -4085 -1432
rect -4131 -2220 -4085 -2208
rect -3973 -1432 -3927 -1420
rect -3973 -2208 -3967 -1432
rect -3933 -2208 -3927 -1432
rect -3973 -2220 -3927 -2208
rect -3815 -1432 -3769 -1420
rect -3815 -2208 -3809 -1432
rect -3775 -2208 -3769 -1432
rect -3815 -2220 -3769 -2208
rect -3657 -1432 -3611 -1420
rect -3657 -2208 -3651 -1432
rect -3617 -2208 -3611 -1432
rect -3657 -2220 -3611 -2208
rect -3499 -1432 -3453 -1420
rect -3499 -2208 -3493 -1432
rect -3459 -2208 -3453 -1432
rect -3499 -2220 -3453 -2208
rect -3341 -1432 -3295 -1420
rect -3341 -2208 -3335 -1432
rect -3301 -2208 -3295 -1432
rect -3341 -2220 -3295 -2208
rect -3183 -1432 -3137 -1420
rect -3183 -2208 -3177 -1432
rect -3143 -2208 -3137 -1432
rect -3183 -2220 -3137 -2208
rect -3025 -1432 -2979 -1420
rect -3025 -2208 -3019 -1432
rect -2985 -2208 -2979 -1432
rect -3025 -2220 -2979 -2208
rect -2867 -1432 -2821 -1420
rect -2867 -2208 -2861 -1432
rect -2827 -2208 -2821 -1432
rect -2867 -2220 -2821 -2208
rect -2709 -1432 -2663 -1420
rect -2709 -2208 -2703 -1432
rect -2669 -2208 -2663 -1432
rect -2709 -2220 -2663 -2208
rect -2551 -1432 -2505 -1420
rect -2551 -2208 -2545 -1432
rect -2511 -2208 -2505 -1432
rect -2551 -2220 -2505 -2208
rect -2393 -1432 -2347 -1420
rect -2393 -2208 -2387 -1432
rect -2353 -2208 -2347 -1432
rect -2393 -2220 -2347 -2208
rect -2235 -1432 -2189 -1420
rect -2235 -2208 -2229 -1432
rect -2195 -2208 -2189 -1432
rect -2235 -2220 -2189 -2208
rect -2077 -1432 -2031 -1420
rect -2077 -2208 -2071 -1432
rect -2037 -2208 -2031 -1432
rect -2077 -2220 -2031 -2208
rect -1919 -1432 -1873 -1420
rect -1919 -2208 -1913 -1432
rect -1879 -2208 -1873 -1432
rect -1919 -2220 -1873 -2208
rect -1761 -1432 -1715 -1420
rect -1761 -2208 -1755 -1432
rect -1721 -2208 -1715 -1432
rect -1761 -2220 -1715 -2208
rect -1603 -1432 -1557 -1420
rect -1603 -2208 -1597 -1432
rect -1563 -2208 -1557 -1432
rect -1603 -2220 -1557 -2208
rect -1445 -1432 -1399 -1420
rect -1445 -2208 -1439 -1432
rect -1405 -2208 -1399 -1432
rect -1445 -2220 -1399 -2208
rect -1287 -1432 -1241 -1420
rect -1287 -2208 -1281 -1432
rect -1247 -2208 -1241 -1432
rect -1287 -2220 -1241 -2208
rect -1129 -1432 -1083 -1420
rect -1129 -2208 -1123 -1432
rect -1089 -2208 -1083 -1432
rect -1129 -2220 -1083 -2208
rect -971 -1432 -925 -1420
rect -971 -2208 -965 -1432
rect -931 -2208 -925 -1432
rect -971 -2220 -925 -2208
rect -813 -1432 -767 -1420
rect -813 -2208 -807 -1432
rect -773 -2208 -767 -1432
rect -813 -2220 -767 -2208
rect -655 -1432 -609 -1420
rect -655 -2208 -649 -1432
rect -615 -2208 -609 -1432
rect -655 -2220 -609 -2208
rect -497 -1432 -451 -1420
rect -497 -2208 -491 -1432
rect -457 -2208 -451 -1432
rect -497 -2220 -451 -2208
rect -339 -1432 -293 -1420
rect -339 -2208 -333 -1432
rect -299 -2208 -293 -1432
rect -339 -2220 -293 -2208
rect -181 -1432 -135 -1420
rect -181 -2208 -175 -1432
rect -141 -2208 -135 -1432
rect -181 -2220 -135 -2208
rect -23 -1432 23 -1420
rect -23 -2208 -17 -1432
rect 17 -2208 23 -1432
rect -23 -2220 23 -2208
rect 135 -1432 181 -1420
rect 135 -2208 141 -1432
rect 175 -2208 181 -1432
rect 135 -2220 181 -2208
rect 293 -1432 339 -1420
rect 293 -2208 299 -1432
rect 333 -2208 339 -1432
rect 293 -2220 339 -2208
rect 451 -1432 497 -1420
rect 451 -2208 457 -1432
rect 491 -2208 497 -1432
rect 451 -2220 497 -2208
rect 609 -1432 655 -1420
rect 609 -2208 615 -1432
rect 649 -2208 655 -1432
rect 609 -2220 655 -2208
rect 767 -1432 813 -1420
rect 767 -2208 773 -1432
rect 807 -2208 813 -1432
rect 767 -2220 813 -2208
rect 925 -1432 971 -1420
rect 925 -2208 931 -1432
rect 965 -2208 971 -1432
rect 925 -2220 971 -2208
rect 1083 -1432 1129 -1420
rect 1083 -2208 1089 -1432
rect 1123 -2208 1129 -1432
rect 1083 -2220 1129 -2208
rect 1241 -1432 1287 -1420
rect 1241 -2208 1247 -1432
rect 1281 -2208 1287 -1432
rect 1241 -2220 1287 -2208
rect 1399 -1432 1445 -1420
rect 1399 -2208 1405 -1432
rect 1439 -2208 1445 -1432
rect 1399 -2220 1445 -2208
rect 1557 -1432 1603 -1420
rect 1557 -2208 1563 -1432
rect 1597 -2208 1603 -1432
rect 1557 -2220 1603 -2208
rect 1715 -1432 1761 -1420
rect 1715 -2208 1721 -1432
rect 1755 -2208 1761 -1432
rect 1715 -2220 1761 -2208
rect 1873 -1432 1919 -1420
rect 1873 -2208 1879 -1432
rect 1913 -2208 1919 -1432
rect 1873 -2220 1919 -2208
rect 2031 -1432 2077 -1420
rect 2031 -2208 2037 -1432
rect 2071 -2208 2077 -1432
rect 2031 -2220 2077 -2208
rect 2189 -1432 2235 -1420
rect 2189 -2208 2195 -1432
rect 2229 -2208 2235 -1432
rect 2189 -2220 2235 -2208
rect 2347 -1432 2393 -1420
rect 2347 -2208 2353 -1432
rect 2387 -2208 2393 -1432
rect 2347 -2220 2393 -2208
rect 2505 -1432 2551 -1420
rect 2505 -2208 2511 -1432
rect 2545 -2208 2551 -1432
rect 2505 -2220 2551 -2208
rect 2663 -1432 2709 -1420
rect 2663 -2208 2669 -1432
rect 2703 -2208 2709 -1432
rect 2663 -2220 2709 -2208
rect 2821 -1432 2867 -1420
rect 2821 -2208 2827 -1432
rect 2861 -2208 2867 -1432
rect 2821 -2220 2867 -2208
rect 2979 -1432 3025 -1420
rect 2979 -2208 2985 -1432
rect 3019 -2208 3025 -1432
rect 2979 -2220 3025 -2208
rect 3137 -1432 3183 -1420
rect 3137 -2208 3143 -1432
rect 3177 -2208 3183 -1432
rect 3137 -2220 3183 -2208
rect 3295 -1432 3341 -1420
rect 3295 -2208 3301 -1432
rect 3335 -2208 3341 -1432
rect 3295 -2220 3341 -2208
rect 3453 -1432 3499 -1420
rect 3453 -2208 3459 -1432
rect 3493 -2208 3499 -1432
rect 3453 -2220 3499 -2208
rect 3611 -1432 3657 -1420
rect 3611 -2208 3617 -1432
rect 3651 -2208 3657 -1432
rect 3611 -2220 3657 -2208
rect 3769 -1432 3815 -1420
rect 3769 -2208 3775 -1432
rect 3809 -2208 3815 -1432
rect 3769 -2220 3815 -2208
rect 3927 -1432 3973 -1420
rect 3927 -2208 3933 -1432
rect 3967 -2208 3973 -1432
rect 3927 -2220 3973 -2208
rect 4085 -1432 4131 -1420
rect 4085 -2208 4091 -1432
rect 4125 -2208 4131 -1432
rect 4085 -2220 4131 -2208
rect 4243 -1432 4289 -1420
rect 4243 -2208 4249 -1432
rect 4283 -2208 4289 -1432
rect 4243 -2220 4289 -2208
rect 4401 -1432 4447 -1420
rect 4401 -2208 4407 -1432
rect 4441 -2208 4447 -1432
rect 4401 -2220 4447 -2208
rect 4559 -1432 4605 -1420
rect 4559 -2208 4565 -1432
rect 4599 -2208 4605 -1432
rect 4559 -2220 4605 -2208
rect 4717 -1432 4763 -1420
rect 4717 -2208 4723 -1432
rect 4757 -2208 4763 -1432
rect 4717 -2220 4763 -2208
rect 4875 -1432 4921 -1420
rect 4875 -2208 4881 -1432
rect 4915 -2208 4921 -1432
rect 4875 -2220 4921 -2208
rect 5033 -1432 5079 -1420
rect 5033 -2208 5039 -1432
rect 5073 -2208 5079 -1432
rect 5033 -2220 5079 -2208
rect 5191 -1432 5237 -1420
rect 5191 -2208 5197 -1432
rect 5231 -2208 5237 -1432
rect 5191 -2220 5237 -2208
rect 5349 -1432 5395 -1420
rect 5349 -2208 5355 -1432
rect 5389 -2208 5395 -1432
rect 5349 -2220 5395 -2208
rect 5507 -1432 5553 -1420
rect 5507 -2208 5513 -1432
rect 5547 -2208 5553 -1432
rect 5507 -2220 5553 -2208
rect 5665 -1432 5711 -1420
rect 5665 -2208 5671 -1432
rect 5705 -2208 5711 -1432
rect 5665 -2220 5711 -2208
rect 5823 -1432 5869 -1420
rect 5823 -2208 5829 -1432
rect 5863 -2208 5869 -1432
rect 5823 -2220 5869 -2208
rect 5981 -1432 6027 -1420
rect 5981 -2208 5987 -1432
rect 6021 -2208 6027 -1432
rect 5981 -2220 6027 -2208
rect 6139 -1432 6185 -1420
rect 6139 -2208 6145 -1432
rect 6179 -2208 6185 -1432
rect 6139 -2220 6185 -2208
rect 6297 -1432 6343 -1420
rect 6297 -2208 6303 -1432
rect 6337 -2208 6343 -1432
rect 6297 -2220 6343 -2208
rect -6287 -2258 -6195 -2252
rect -6287 -2292 -6275 -2258
rect -6207 -2292 -6195 -2258
rect -6287 -2298 -6195 -2292
rect -6129 -2258 -6037 -2252
rect -6129 -2292 -6117 -2258
rect -6049 -2292 -6037 -2258
rect -6129 -2298 -6037 -2292
rect -5971 -2258 -5879 -2252
rect -5971 -2292 -5959 -2258
rect -5891 -2292 -5879 -2258
rect -5971 -2298 -5879 -2292
rect -5813 -2258 -5721 -2252
rect -5813 -2292 -5801 -2258
rect -5733 -2292 -5721 -2258
rect -5813 -2298 -5721 -2292
rect -5655 -2258 -5563 -2252
rect -5655 -2292 -5643 -2258
rect -5575 -2292 -5563 -2258
rect -5655 -2298 -5563 -2292
rect -5497 -2258 -5405 -2252
rect -5497 -2292 -5485 -2258
rect -5417 -2292 -5405 -2258
rect -5497 -2298 -5405 -2292
rect -5339 -2258 -5247 -2252
rect -5339 -2292 -5327 -2258
rect -5259 -2292 -5247 -2258
rect -5339 -2298 -5247 -2292
rect -5181 -2258 -5089 -2252
rect -5181 -2292 -5169 -2258
rect -5101 -2292 -5089 -2258
rect -5181 -2298 -5089 -2292
rect -5023 -2258 -4931 -2252
rect -5023 -2292 -5011 -2258
rect -4943 -2292 -4931 -2258
rect -5023 -2298 -4931 -2292
rect -4865 -2258 -4773 -2252
rect -4865 -2292 -4853 -2258
rect -4785 -2292 -4773 -2258
rect -4865 -2298 -4773 -2292
rect -4707 -2258 -4615 -2252
rect -4707 -2292 -4695 -2258
rect -4627 -2292 -4615 -2258
rect -4707 -2298 -4615 -2292
rect -4549 -2258 -4457 -2252
rect -4549 -2292 -4537 -2258
rect -4469 -2292 -4457 -2258
rect -4549 -2298 -4457 -2292
rect -4391 -2258 -4299 -2252
rect -4391 -2292 -4379 -2258
rect -4311 -2292 -4299 -2258
rect -4391 -2298 -4299 -2292
rect -4233 -2258 -4141 -2252
rect -4233 -2292 -4221 -2258
rect -4153 -2292 -4141 -2258
rect -4233 -2298 -4141 -2292
rect -4075 -2258 -3983 -2252
rect -4075 -2292 -4063 -2258
rect -3995 -2292 -3983 -2258
rect -4075 -2298 -3983 -2292
rect -3917 -2258 -3825 -2252
rect -3917 -2292 -3905 -2258
rect -3837 -2292 -3825 -2258
rect -3917 -2298 -3825 -2292
rect -3759 -2258 -3667 -2252
rect -3759 -2292 -3747 -2258
rect -3679 -2292 -3667 -2258
rect -3759 -2298 -3667 -2292
rect -3601 -2258 -3509 -2252
rect -3601 -2292 -3589 -2258
rect -3521 -2292 -3509 -2258
rect -3601 -2298 -3509 -2292
rect -3443 -2258 -3351 -2252
rect -3443 -2292 -3431 -2258
rect -3363 -2292 -3351 -2258
rect -3443 -2298 -3351 -2292
rect -3285 -2258 -3193 -2252
rect -3285 -2292 -3273 -2258
rect -3205 -2292 -3193 -2258
rect -3285 -2298 -3193 -2292
rect -3127 -2258 -3035 -2252
rect -3127 -2292 -3115 -2258
rect -3047 -2292 -3035 -2258
rect -3127 -2298 -3035 -2292
rect -2969 -2258 -2877 -2252
rect -2969 -2292 -2957 -2258
rect -2889 -2292 -2877 -2258
rect -2969 -2298 -2877 -2292
rect -2811 -2258 -2719 -2252
rect -2811 -2292 -2799 -2258
rect -2731 -2292 -2719 -2258
rect -2811 -2298 -2719 -2292
rect -2653 -2258 -2561 -2252
rect -2653 -2292 -2641 -2258
rect -2573 -2292 -2561 -2258
rect -2653 -2298 -2561 -2292
rect -2495 -2258 -2403 -2252
rect -2495 -2292 -2483 -2258
rect -2415 -2292 -2403 -2258
rect -2495 -2298 -2403 -2292
rect -2337 -2258 -2245 -2252
rect -2337 -2292 -2325 -2258
rect -2257 -2292 -2245 -2258
rect -2337 -2298 -2245 -2292
rect -2179 -2258 -2087 -2252
rect -2179 -2292 -2167 -2258
rect -2099 -2292 -2087 -2258
rect -2179 -2298 -2087 -2292
rect -2021 -2258 -1929 -2252
rect -2021 -2292 -2009 -2258
rect -1941 -2292 -1929 -2258
rect -2021 -2298 -1929 -2292
rect -1863 -2258 -1771 -2252
rect -1863 -2292 -1851 -2258
rect -1783 -2292 -1771 -2258
rect -1863 -2298 -1771 -2292
rect -1705 -2258 -1613 -2252
rect -1705 -2292 -1693 -2258
rect -1625 -2292 -1613 -2258
rect -1705 -2298 -1613 -2292
rect -1547 -2258 -1455 -2252
rect -1547 -2292 -1535 -2258
rect -1467 -2292 -1455 -2258
rect -1547 -2298 -1455 -2292
rect -1389 -2258 -1297 -2252
rect -1389 -2292 -1377 -2258
rect -1309 -2292 -1297 -2258
rect -1389 -2298 -1297 -2292
rect -1231 -2258 -1139 -2252
rect -1231 -2292 -1219 -2258
rect -1151 -2292 -1139 -2258
rect -1231 -2298 -1139 -2292
rect -1073 -2258 -981 -2252
rect -1073 -2292 -1061 -2258
rect -993 -2292 -981 -2258
rect -1073 -2298 -981 -2292
rect -915 -2258 -823 -2252
rect -915 -2292 -903 -2258
rect -835 -2292 -823 -2258
rect -915 -2298 -823 -2292
rect -757 -2258 -665 -2252
rect -757 -2292 -745 -2258
rect -677 -2292 -665 -2258
rect -757 -2298 -665 -2292
rect -599 -2258 -507 -2252
rect -599 -2292 -587 -2258
rect -519 -2292 -507 -2258
rect -599 -2298 -507 -2292
rect -441 -2258 -349 -2252
rect -441 -2292 -429 -2258
rect -361 -2292 -349 -2258
rect -441 -2298 -349 -2292
rect -283 -2258 -191 -2252
rect -283 -2292 -271 -2258
rect -203 -2292 -191 -2258
rect -283 -2298 -191 -2292
rect -125 -2258 -33 -2252
rect -125 -2292 -113 -2258
rect -45 -2292 -33 -2258
rect -125 -2298 -33 -2292
rect 33 -2258 125 -2252
rect 33 -2292 45 -2258
rect 113 -2292 125 -2258
rect 33 -2298 125 -2292
rect 191 -2258 283 -2252
rect 191 -2292 203 -2258
rect 271 -2292 283 -2258
rect 191 -2298 283 -2292
rect 349 -2258 441 -2252
rect 349 -2292 361 -2258
rect 429 -2292 441 -2258
rect 349 -2298 441 -2292
rect 507 -2258 599 -2252
rect 507 -2292 519 -2258
rect 587 -2292 599 -2258
rect 507 -2298 599 -2292
rect 665 -2258 757 -2252
rect 665 -2292 677 -2258
rect 745 -2292 757 -2258
rect 665 -2298 757 -2292
rect 823 -2258 915 -2252
rect 823 -2292 835 -2258
rect 903 -2292 915 -2258
rect 823 -2298 915 -2292
rect 981 -2258 1073 -2252
rect 981 -2292 993 -2258
rect 1061 -2292 1073 -2258
rect 981 -2298 1073 -2292
rect 1139 -2258 1231 -2252
rect 1139 -2292 1151 -2258
rect 1219 -2292 1231 -2258
rect 1139 -2298 1231 -2292
rect 1297 -2258 1389 -2252
rect 1297 -2292 1309 -2258
rect 1377 -2292 1389 -2258
rect 1297 -2298 1389 -2292
rect 1455 -2258 1547 -2252
rect 1455 -2292 1467 -2258
rect 1535 -2292 1547 -2258
rect 1455 -2298 1547 -2292
rect 1613 -2258 1705 -2252
rect 1613 -2292 1625 -2258
rect 1693 -2292 1705 -2258
rect 1613 -2298 1705 -2292
rect 1771 -2258 1863 -2252
rect 1771 -2292 1783 -2258
rect 1851 -2292 1863 -2258
rect 1771 -2298 1863 -2292
rect 1929 -2258 2021 -2252
rect 1929 -2292 1941 -2258
rect 2009 -2292 2021 -2258
rect 1929 -2298 2021 -2292
rect 2087 -2258 2179 -2252
rect 2087 -2292 2099 -2258
rect 2167 -2292 2179 -2258
rect 2087 -2298 2179 -2292
rect 2245 -2258 2337 -2252
rect 2245 -2292 2257 -2258
rect 2325 -2292 2337 -2258
rect 2245 -2298 2337 -2292
rect 2403 -2258 2495 -2252
rect 2403 -2292 2415 -2258
rect 2483 -2292 2495 -2258
rect 2403 -2298 2495 -2292
rect 2561 -2258 2653 -2252
rect 2561 -2292 2573 -2258
rect 2641 -2292 2653 -2258
rect 2561 -2298 2653 -2292
rect 2719 -2258 2811 -2252
rect 2719 -2292 2731 -2258
rect 2799 -2292 2811 -2258
rect 2719 -2298 2811 -2292
rect 2877 -2258 2969 -2252
rect 2877 -2292 2889 -2258
rect 2957 -2292 2969 -2258
rect 2877 -2298 2969 -2292
rect 3035 -2258 3127 -2252
rect 3035 -2292 3047 -2258
rect 3115 -2292 3127 -2258
rect 3035 -2298 3127 -2292
rect 3193 -2258 3285 -2252
rect 3193 -2292 3205 -2258
rect 3273 -2292 3285 -2258
rect 3193 -2298 3285 -2292
rect 3351 -2258 3443 -2252
rect 3351 -2292 3363 -2258
rect 3431 -2292 3443 -2258
rect 3351 -2298 3443 -2292
rect 3509 -2258 3601 -2252
rect 3509 -2292 3521 -2258
rect 3589 -2292 3601 -2258
rect 3509 -2298 3601 -2292
rect 3667 -2258 3759 -2252
rect 3667 -2292 3679 -2258
rect 3747 -2292 3759 -2258
rect 3667 -2298 3759 -2292
rect 3825 -2258 3917 -2252
rect 3825 -2292 3837 -2258
rect 3905 -2292 3917 -2258
rect 3825 -2298 3917 -2292
rect 3983 -2258 4075 -2252
rect 3983 -2292 3995 -2258
rect 4063 -2292 4075 -2258
rect 3983 -2298 4075 -2292
rect 4141 -2258 4233 -2252
rect 4141 -2292 4153 -2258
rect 4221 -2292 4233 -2258
rect 4141 -2298 4233 -2292
rect 4299 -2258 4391 -2252
rect 4299 -2292 4311 -2258
rect 4379 -2292 4391 -2258
rect 4299 -2298 4391 -2292
rect 4457 -2258 4549 -2252
rect 4457 -2292 4469 -2258
rect 4537 -2292 4549 -2258
rect 4457 -2298 4549 -2292
rect 4615 -2258 4707 -2252
rect 4615 -2292 4627 -2258
rect 4695 -2292 4707 -2258
rect 4615 -2298 4707 -2292
rect 4773 -2258 4865 -2252
rect 4773 -2292 4785 -2258
rect 4853 -2292 4865 -2258
rect 4773 -2298 4865 -2292
rect 4931 -2258 5023 -2252
rect 4931 -2292 4943 -2258
rect 5011 -2292 5023 -2258
rect 4931 -2298 5023 -2292
rect 5089 -2258 5181 -2252
rect 5089 -2292 5101 -2258
rect 5169 -2292 5181 -2258
rect 5089 -2298 5181 -2292
rect 5247 -2258 5339 -2252
rect 5247 -2292 5259 -2258
rect 5327 -2292 5339 -2258
rect 5247 -2298 5339 -2292
rect 5405 -2258 5497 -2252
rect 5405 -2292 5417 -2258
rect 5485 -2292 5497 -2258
rect 5405 -2298 5497 -2292
rect 5563 -2258 5655 -2252
rect 5563 -2292 5575 -2258
rect 5643 -2292 5655 -2258
rect 5563 -2298 5655 -2292
rect 5721 -2258 5813 -2252
rect 5721 -2292 5733 -2258
rect 5801 -2292 5813 -2258
rect 5721 -2298 5813 -2292
rect 5879 -2258 5971 -2252
rect 5879 -2292 5891 -2258
rect 5959 -2292 5971 -2258
rect 5879 -2298 5971 -2292
rect 6037 -2258 6129 -2252
rect 6037 -2292 6049 -2258
rect 6117 -2292 6129 -2258
rect 6037 -2298 6129 -2292
rect 6195 -2258 6287 -2252
rect 6195 -2292 6207 -2258
rect 6275 -2292 6287 -2258
rect 6195 -2298 6287 -2292
<< properties >>
string FIXED_BBOX -6454 -2413 6454 2413
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.50 m 5 nf 80 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
