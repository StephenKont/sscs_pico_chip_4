magic
tech sky130A
magscale 1 2
timestamp 1667858459
<< viali >>
rect 467844 450395 468039 450429
rect 468206 450395 468402 450429
rect 468844 450395 469039 450429
rect 469206 450395 469402 450429
rect 467748 449775 467782 450333
rect 468054 450185 468192 450219
rect 467958 449985 467992 450123
rect 468090 450021 468156 450087
rect 468254 449985 468288 450123
rect 468464 449775 468498 450333
rect 468748 449775 468782 450333
rect 469054 450185 469192 450219
rect 468958 449985 468992 450123
rect 469090 450021 469156 450087
rect 469254 449985 469288 450123
rect 469464 449775 469498 450333
rect 467844 449679 468402 449713
rect 468844 449679 469402 449713
rect 334420 389741 334615 389775
rect 334782 389741 334978 389775
rect 335420 389741 335615 389775
rect 335782 389741 335978 389775
rect 334324 389121 334358 389679
rect 334630 389531 334768 389565
rect 334534 389331 334568 389469
rect 334830 389331 334864 389469
rect 335040 389121 335074 389679
rect 335324 389121 335358 389679
rect 335630 389531 335768 389565
rect 335534 389331 335568 389469
rect 335830 389331 335864 389469
rect 336040 389121 336074 389679
rect 334420 389025 334978 389059
rect 335420 389025 335978 389059
<< metal1 >>
rect 351259 697923 404827 699695
rect 406599 697923 406605 699695
rect 145394 681965 165394 682901
rect 145394 674731 146520 681965
rect 164088 674731 165394 681965
rect 145394 567969 165394 674731
rect 351259 610221 353031 697923
rect 529662 696917 530093 696928
rect 529662 696526 529691 696917
rect 530082 696526 533502 696917
rect 529662 696509 530093 696526
rect 418923 692927 531009 693157
rect 418923 690516 419153 692927
rect 418001 690286 419153 690516
rect 530779 685003 531009 692927
rect 533111 691809 533502 696526
rect 533111 691418 535568 691809
rect 540110 687288 540426 687322
rect 540110 687119 540137 687288
rect 540399 687119 540426 687288
rect 540110 687092 540426 687119
rect 540143 685003 540373 687092
rect 530779 684773 540373 685003
rect 540143 684600 540373 684773
rect 540143 684370 571624 684600
rect 442918 679662 462918 680730
rect 442918 669616 443952 679662
rect 462134 669616 462918 679662
rect 442918 613648 462918 669616
rect 442918 599950 444062 613648
rect 461834 599950 462918 613648
rect 442918 598730 462918 599950
rect 145394 556095 146784 567969
rect 164076 556095 165394 567969
rect 145394 553901 165394 556095
rect 145398 511617 165398 512903
rect 145398 498073 146694 511617
rect 163458 498073 165398 511617
rect 145398 409147 165398 498073
rect 468092 460164 468156 460170
rect 467736 450441 468045 450442
rect 467735 450429 468045 450441
rect 467735 450395 467844 450429
rect 468039 450395 468045 450429
rect 467735 450383 468045 450395
rect 467735 450333 467794 450383
rect 467735 449775 467748 450333
rect 467782 449775 467794 450333
rect 468092 450231 468156 460100
rect 469092 458678 469156 458684
rect 468200 450429 468510 450442
rect 468736 450441 469045 450442
rect 468200 450395 468206 450429
rect 468402 450395 468510 450429
rect 468200 450383 468510 450395
rect 468452 450333 468510 450383
rect 467946 450219 468300 450231
rect 467946 450185 468054 450219
rect 468192 450185 468300 450219
rect 467946 450173 468300 450185
rect 467946 450123 468004 450173
rect 467946 449985 467958 450123
rect 467992 449985 468004 450123
rect 468242 450123 468300 450173
rect 467946 449877 468004 449985
rect 468078 450087 468168 450099
rect 468078 450021 468090 450087
rect 468156 450021 468168 450087
rect 467735 449725 467794 449775
rect 468078 449725 468168 450021
rect 468242 449985 468254 450123
rect 468288 449985 468300 450123
rect 468242 449877 468300 449985
rect 468452 449775 468464 450333
rect 468498 449775 468510 450333
rect 468452 449725 468510 449775
rect 467735 449713 468510 449725
rect 467735 449679 467844 449713
rect 468402 449679 468510 449713
rect 467735 449667 468510 449679
rect 467735 449521 467794 449667
rect 468452 449521 468510 449667
rect 468735 450429 469045 450441
rect 468735 450395 468844 450429
rect 469039 450395 469045 450429
rect 468735 450383 469045 450395
rect 468735 450333 468794 450383
rect 468735 449775 468748 450333
rect 468782 449775 468794 450333
rect 469092 450231 469156 458614
rect 469200 450429 469510 450442
rect 469200 450395 469206 450429
rect 469402 450395 469510 450429
rect 469200 450383 469510 450395
rect 469452 450333 469510 450383
rect 468946 450219 469300 450231
rect 468946 450185 469054 450219
rect 469192 450185 469300 450219
rect 468946 450173 469300 450185
rect 468946 450123 469004 450173
rect 468946 449985 468958 450123
rect 468992 449985 469004 450123
rect 469242 450123 469300 450173
rect 468946 449877 469004 449985
rect 469078 450087 469168 450099
rect 469078 450021 469090 450087
rect 469156 450021 469168 450087
rect 468735 449725 468794 449775
rect 469078 449725 469168 450021
rect 469242 449985 469254 450123
rect 469288 449985 469300 450123
rect 469242 449877 469300 449985
rect 469452 449775 469464 450333
rect 469498 449775 469510 450333
rect 469452 449725 469510 449775
rect 468735 449713 469510 449725
rect 468735 449679 468844 449713
rect 469402 449679 469510 449713
rect 468735 449667 469510 449679
rect 468735 449521 468794 449667
rect 469452 449521 469510 449667
rect 467580 449507 469674 449521
rect 467580 449422 467592 449507
rect 469659 449422 469674 449507
rect 467580 449411 469674 449422
rect 145398 401839 146500 409147
rect 164068 401839 165398 409147
rect 145398 400903 165398 401839
rect 335657 390802 335741 390811
rect 335657 390738 335668 390802
rect 335732 390738 335741 390802
rect 335657 390728 335741 390738
rect 334650 390146 334758 390164
rect 334650 390082 334668 390146
rect 334732 390082 334758 390146
rect 334650 390066 334758 390082
rect 334312 389787 334621 389788
rect 334311 389775 334621 389787
rect 334311 389741 334420 389775
rect 334615 389741 334621 389775
rect 334311 389729 334621 389741
rect 334311 389679 334370 389729
rect 334311 389121 334324 389679
rect 334358 389121 334370 389679
rect 334668 389577 334732 390066
rect 334776 389775 335086 389788
rect 335312 389787 335621 389788
rect 334776 389741 334782 389775
rect 334978 389741 335086 389775
rect 334776 389729 335086 389741
rect 335028 389679 335086 389729
rect 334522 389565 334876 389577
rect 334522 389531 334630 389565
rect 334768 389531 334876 389565
rect 334522 389519 334876 389531
rect 334522 389469 334580 389519
rect 334522 389331 334534 389469
rect 334568 389331 334580 389469
rect 334818 389469 334876 389519
rect 334522 389223 334580 389331
rect 334311 389071 334370 389121
rect 334654 389071 334744 389445
rect 334818 389331 334830 389469
rect 334864 389331 334876 389469
rect 334818 389223 334876 389331
rect 335028 389121 335040 389679
rect 335074 389121 335086 389679
rect 335028 389071 335086 389121
rect 334311 389059 335086 389071
rect 334311 389025 334420 389059
rect 334978 389025 335086 389059
rect 334311 389013 335086 389025
rect 334311 388853 334370 389013
rect 335028 388853 335086 389013
rect 335311 389775 335621 389787
rect 335311 389741 335420 389775
rect 335615 389741 335621 389775
rect 335311 389729 335621 389741
rect 335311 389679 335370 389729
rect 335311 389121 335324 389679
rect 335358 389121 335370 389679
rect 335668 389577 335732 390728
rect 335776 389775 336086 389788
rect 335776 389741 335782 389775
rect 335978 389741 336086 389775
rect 335776 389729 336086 389741
rect 336028 389679 336086 389729
rect 335522 389565 335876 389577
rect 335522 389531 335630 389565
rect 335768 389531 335876 389565
rect 335522 389519 335876 389531
rect 335522 389469 335580 389519
rect 335522 389331 335534 389469
rect 335568 389331 335580 389469
rect 335818 389469 335876 389519
rect 335522 389223 335580 389331
rect 335311 389071 335370 389121
rect 335654 389071 335744 389445
rect 335818 389331 335830 389469
rect 335864 389331 335876 389469
rect 335818 389223 335876 389331
rect 336028 389121 336040 389679
rect 336074 389121 336086 389679
rect 336028 389071 336086 389121
rect 335311 389059 336086 389071
rect 335311 389025 335420 389059
rect 335978 389025 336086 389059
rect 335311 389013 336086 389025
rect 335311 388853 335370 389013
rect 336028 388853 336086 389013
rect 333727 388772 336528 388853
rect 333727 387884 333824 388772
rect 336416 387884 336528 388772
rect 333727 387811 336528 387884
<< via1 >>
rect 404827 697923 406599 699695
rect 146520 674731 164088 681965
rect 529691 696526 530082 696917
rect 540137 687119 540399 687288
rect 443952 669616 462134 679662
rect 444062 599950 461834 613648
rect 146784 556095 164076 567969
rect 146694 498073 163458 511617
rect 468092 460100 468156 460164
rect 469092 458614 469156 458678
rect 467592 449422 469659 449507
rect 146500 401839 164068 409147
rect 335668 390738 335732 390802
rect 334668 390082 334732 390146
rect 333824 387884 336416 388772
<< metal2 >>
rect 404827 699695 406599 699701
rect 404818 697923 404827 699695
rect 406599 697923 406608 699695
rect 404827 697917 406599 697923
rect 529662 696917 530093 696928
rect 529662 696526 529691 696917
rect 530082 696526 530093 696917
rect 529662 696509 530093 696526
rect 326218 693564 337501 693970
rect 326218 692489 326803 693564
rect 327878 693559 337501 693564
rect 327878 692494 335984 693559
rect 337049 692494 337501 693559
rect 327878 692489 337501 692494
rect 326218 691947 337501 692489
rect 434817 687328 525966 688544
rect 145394 681965 165394 682901
rect 145394 674731 146520 681965
rect 164088 674731 165394 681965
rect 416733 680130 417949 680139
rect 416733 676381 417949 678914
rect 434817 676381 436033 687328
rect 524750 682605 525966 687328
rect 540110 687288 540426 687322
rect 540110 687119 540137 687288
rect 540399 687119 540426 687288
rect 540110 687092 540426 687119
rect 524750 681389 571624 682605
rect 416733 675165 436033 676381
rect 442918 679662 462918 680730
rect 145394 567969 165394 674731
rect 442918 669616 443952 679662
rect 462134 669616 462918 679662
rect 442918 613648 462918 669616
rect 442918 599950 444062 613648
rect 461834 599950 462918 613648
rect 442918 598730 462918 599950
rect 145394 556095 146784 567969
rect 164076 556095 165394 567969
rect 145394 553901 165394 556095
rect 145398 511617 165398 512903
rect 145398 498073 146694 511617
rect 163458 498073 165398 511617
rect 145398 409147 165398 498073
rect 468083 460100 468092 460164
rect 468156 460100 468165 460164
rect 469083 458614 469092 458678
rect 469156 458614 469165 458678
rect 467580 449507 469674 449521
rect 467580 449422 467592 449507
rect 469659 449422 469674 449507
rect 467580 449411 469674 449422
rect 145398 401839 146500 409147
rect 164068 401839 165398 409147
rect 315391 430218 315511 430227
rect 315391 404023 315407 430218
rect 315496 404023 315511 430218
rect 315391 404007 315511 404023
rect 145398 400903 165398 401839
rect 335657 390802 335741 390811
rect 335657 390738 335668 390802
rect 335732 390738 335741 390802
rect 335657 390728 335741 390738
rect 334650 390146 334758 390164
rect 334650 390082 334668 390146
rect 334732 390082 334758 390146
rect 334650 390066 334758 390082
rect 333727 388772 336528 388853
rect 333727 387884 333824 388772
rect 336416 387884 336528 388772
rect 333727 387811 336528 387884
<< via2 >>
rect 550609 700259 558926 701830
rect 404827 697923 406599 699695
rect 529691 696526 530082 696917
rect 326803 692489 327878 693564
rect 335984 692494 337049 693559
rect 551759 687343 558970 687415
rect 146520 674731 164088 681965
rect 416733 678914 417949 680130
rect 550549 687127 558970 687343
rect 550549 686454 551847 687127
rect 443952 669616 462134 679662
rect 444062 599950 461834 613648
rect 146784 556095 164076 567969
rect 146694 498073 163458 511617
rect 468092 460100 468156 460164
rect 469092 458614 469156 458678
rect 467592 449422 469659 449507
rect 146500 401839 164068 409147
rect 315407 404023 315496 430218
rect 335668 390738 335732 390802
rect 334668 390082 334732 390146
rect 333824 387884 336416 388772
<< metal3 >>
rect 550498 701830 564228 703732
rect 550498 700259 550609 701830
rect 558926 700259 564228 701830
rect 550498 700176 564228 700259
rect 68194 693228 73194 697520
rect 120194 695306 196134 700140
rect 68194 688228 182550 693228
rect 35194 682901 163994 685390
rect 177550 682901 182550 688228
rect 191134 692480 196134 695306
rect 326798 693564 327883 693569
rect 319829 692489 319835 693564
rect 320910 692489 326803 693564
rect 327878 692489 327883 693564
rect 326798 692484 327883 692489
rect 191134 687480 212060 692480
rect 207060 683876 212060 687480
rect 35194 681965 165394 682901
rect 35194 680390 146520 681965
rect 37396 680389 146520 680390
rect 145394 674731 146520 680389
rect 164088 674731 165394 681965
rect 145394 672901 165394 674731
rect 177396 681741 193396 682901
rect 177396 673993 178294 681741
rect 192634 673993 193396 681741
rect 207060 678876 310182 683876
rect 207060 678875 301396 678876
rect 177396 671901 193396 673993
rect 177396 655901 301396 671901
rect 37396 638901 284396 654901
rect 37396 427901 53396 638901
rect 54396 621901 267396 637901
rect 54396 444901 70396 621901
rect 71396 604901 250396 620901
rect 71396 461901 87396 604901
rect 88396 587901 233396 603901
rect 88396 478901 104396 587901
rect 105396 570901 216396 586901
rect 105396 495901 121396 570901
rect 145394 567969 165394 569901
rect 145394 556095 146784 567969
rect 164076 556095 165394 567969
rect 145394 553901 165394 556095
rect 200396 512901 216396 570901
rect 145398 511617 216396 512901
rect 145398 498073 146694 511617
rect 163458 498073 216396 511617
rect 145398 496787 216396 498073
rect 217396 495901 233396 587901
rect 105396 479901 233396 495901
rect 234396 478901 250396 604901
rect 88396 462901 250396 478901
rect 251396 461901 267396 621901
rect 71396 445901 267396 461901
rect 268396 444901 284396 638901
rect 54396 428901 284396 444901
rect 285396 427901 301396 655901
rect 305182 614574 310182 678876
rect 329491 669335 333977 700140
rect 404822 699695 406604 699700
rect 415342 699695 417114 700140
rect 404822 697923 404827 699695
rect 406599 697926 417114 699695
rect 406599 697923 408680 697926
rect 404822 697918 406604 697923
rect 465394 695162 470394 700140
rect 335979 693559 409017 693564
rect 335979 692494 335984 693559
rect 337049 692494 409017 693559
rect 335979 692489 409017 692494
rect 407942 678700 409017 692489
rect 465394 692349 507525 695162
rect 509588 694218 510140 700140
rect 525390 694218 525836 700140
rect 529662 696922 530093 696928
rect 529662 696521 529686 696922
rect 530077 696917 530093 696922
rect 530082 696526 530093 696917
rect 530077 696521 530093 696526
rect 529662 696509 530093 696521
rect 509588 693836 525836 694218
rect 465394 690162 526363 692349
rect 523478 686995 526363 690162
rect 550247 687533 552095 687538
rect 550247 687415 559057 687533
rect 550247 687343 551759 687415
rect 550247 686995 550549 687343
rect 558970 687127 559057 687415
rect 523478 686454 550549 686995
rect 551847 686454 559057 687127
rect 523478 685110 559057 686454
rect 416733 680135 417949 680886
rect 416728 680130 417954 680135
rect 416728 678914 416733 680130
rect 417949 678914 417954 680130
rect 416728 678909 417954 678914
rect 442918 679662 462918 680730
rect 407942 678617 422717 678700
rect 407942 677625 430204 678617
rect 442918 669616 443952 679662
rect 462134 669616 462918 679662
rect 472300 680688 571624 682984
rect 472300 676484 472834 680688
rect 491834 677984 571624 680688
rect 491834 676484 492300 677984
rect 472300 675984 492300 676484
rect 442918 668730 462918 669616
rect 442918 664966 567918 665730
rect 442918 650540 443558 664966
rect 462290 650540 567918 664966
rect 442918 649730 567918 650540
rect 365918 632730 550918 648730
rect 305182 613572 334874 614574
rect 365918 483730 381918 632730
rect 382918 615730 533918 631730
rect 382918 500730 398918 615730
rect 399918 613648 462918 614730
rect 399918 599950 444062 613648
rect 461834 599950 462918 613648
rect 399918 598730 462918 599950
rect 399918 517730 415918 598730
rect 517918 517730 533918 615730
rect 399918 501730 533918 517730
rect 534918 500730 550918 632730
rect 382918 484730 550918 500730
rect 551918 483730 567918 649730
rect 365918 467730 567918 483730
rect 359782 460164 571624 460259
rect 359782 460100 468092 460164
rect 468156 460100 571624 460164
rect 359782 460029 571624 460100
rect 37396 411901 301396 427901
rect 315391 430218 315511 430227
rect 145398 409147 165398 410903
rect 145398 403732 146500 409147
rect 35194 401839 146500 403732
rect 164068 401839 165398 409147
rect 315391 404023 315407 430218
rect 315496 404023 315511 430218
rect 315391 404007 315511 404023
rect 35194 400903 165398 401839
rect 35194 398732 164798 400903
rect 359782 393971 360012 460029
rect 345229 393741 360012 393971
rect 364943 458678 571624 458843
rect 364943 458614 469092 458678
rect 469156 458614 571624 458678
rect 364943 458415 571624 458614
rect 335668 391085 335732 391091
rect 335668 390811 335732 391021
rect 345229 390883 345459 393741
rect 364943 393188 365371 458415
rect 467580 449507 469674 449521
rect 467580 449422 467592 449507
rect 469659 449422 469674 449507
rect 467580 449411 469674 449422
rect 359664 392760 365371 393188
rect 335657 390802 335741 390811
rect 335657 390738 335668 390802
rect 335732 390738 335741 390802
rect 335657 390728 335741 390738
rect 334650 390151 334758 390164
rect 334650 390077 334663 390151
rect 334737 390077 334758 390151
rect 334650 390066 334758 390077
rect 333727 388772 336528 388853
rect 333727 387884 333824 388772
rect 336416 387884 336528 388772
rect 333727 387811 336528 387884
<< rmetal3 >>
rect 67397 697520 73795 700140
<< via3 >>
rect 319835 692489 320910 693564
rect 146520 674731 164088 681965
rect 178294 673993 192634 681741
rect 146784 556095 164076 567969
rect 510140 694218 525390 700140
rect 529686 696917 530077 696922
rect 529686 696526 529691 696917
rect 529691 696526 530077 696917
rect 529686 696521 530077 696526
rect 443952 669616 462134 679662
rect 472834 676484 491834 680688
rect 329310 625656 329890 666846
rect 443558 650540 462290 664966
rect 327010 615420 327590 625656
rect 146500 401839 164068 409147
rect 315407 404023 315496 430218
rect 335668 391021 335732 391085
rect 467592 449422 469659 449507
rect 334663 390146 334737 390151
rect 334663 390082 334668 390146
rect 334668 390082 334732 390146
rect 334732 390082 334737 390146
rect 334663 390077 334737 390082
rect 333824 387884 336416 388772
<< metal4 >>
rect 509482 700140 525794 700828
rect 217076 694329 313018 700140
rect 217076 694064 326008 694329
rect 303443 693564 326008 694064
rect 303443 692489 319835 693564
rect 320910 692489 326008 693564
rect 303443 685915 326008 692489
rect 145394 681965 165394 682901
rect 145394 674731 146520 681965
rect 164088 674731 165394 681965
rect 145394 672901 165394 674731
rect 177396 681741 193396 682901
rect 177396 673993 178294 681741
rect 192634 673993 193396 681741
rect 177396 672901 193396 673993
rect 37396 655903 301396 671903
rect 318008 668449 326008 685915
rect 329491 680766 333977 700140
rect 344882 694218 510140 700140
rect 525390 696917 525836 700140
rect 529662 696922 530093 696928
rect 529662 696917 529686 696922
rect 525390 696526 529686 696917
rect 525390 694218 525836 696526
rect 529662 696521 529686 696526
rect 530077 696521 530093 696922
rect 529662 696509 530093 696521
rect 344882 694016 525836 694218
rect 329491 669335 333996 680766
rect 344882 679466 352882 694016
rect 509588 693836 525836 694016
rect 419347 680730 454676 683321
rect 419347 680128 462918 680730
rect 344618 671466 352882 679466
rect 318008 667405 326803 668449
rect 318008 666882 329224 667405
rect 318008 666856 329488 666882
rect 318008 666846 329900 666856
rect 37396 427903 53396 655903
rect 54394 638901 284394 654901
rect 54394 444901 70394 638901
rect 71394 621901 267394 637901
rect 71394 461901 87394 621901
rect 88394 604901 250394 620901
rect 88394 478901 104394 604901
rect 105394 587901 233394 604017
rect 105394 495901 121394 587901
rect 122394 567969 165394 569901
rect 122394 556095 146784 567969
rect 164076 556095 165394 567969
rect 122394 553901 165394 556095
rect 122394 512901 138394 553901
rect 217394 512901 233394 587901
rect 122394 496901 233394 512901
rect 234394 495901 250394 604901
rect 105394 479901 250394 495901
rect 251394 478901 267394 621901
rect 88394 462901 267394 478901
rect 268394 461901 284394 638901
rect 71394 445901 284394 461901
rect 285394 444901 301394 655903
rect 318008 641449 329310 666846
rect 320810 625656 329310 641449
rect 329890 625656 329900 666846
rect 333349 625826 333996 669335
rect 344882 650788 352882 671466
rect 442918 679662 462918 680128
rect 442918 669616 443952 679662
rect 462134 669616 462918 679662
rect 472300 680688 492300 680984
rect 472300 676484 472834 680688
rect 491834 676484 492300 680688
rect 472300 675984 492300 676484
rect 442918 668730 462918 669616
rect 365918 664966 462918 665730
rect 365918 650540 443558 664966
rect 462290 650540 462918 664966
rect 365918 649730 462918 650540
rect 320810 625646 327010 625656
rect 327000 615420 327010 625646
rect 327590 625646 329900 625656
rect 327590 615420 327600 625646
rect 327000 615410 327600 615420
rect 355680 594766 356922 618535
rect 345203 593524 356922 594766
rect 345203 453097 346445 593524
rect 365918 483730 381918 649730
rect 382918 632730 567918 648730
rect 382918 500730 398918 632730
rect 399918 615730 550918 631730
rect 399918 517730 415918 615730
rect 470918 613524 533918 614730
rect 470918 599798 472272 613524
rect 489906 599798 533918 613524
rect 470918 598730 533918 599798
rect 517918 517730 533918 598730
rect 399918 501730 533918 517730
rect 534918 500730 550918 615730
rect 382918 484730 550918 500730
rect 551918 483730 567918 632730
rect 365918 467730 567918 483730
rect 350636 460921 385103 460945
rect 350636 455969 350660 460921
rect 355612 456299 385103 460921
rect 355612 455969 380103 456299
rect 350636 455945 380103 455969
rect 345203 451855 364263 453097
rect 363221 449507 364263 451855
rect 467580 449507 469674 449521
rect 363221 449422 467592 449507
rect 469659 449422 484266 449507
rect 363221 448557 484266 449422
rect 363841 445744 484266 448557
rect 54394 428901 301394 444901
rect 315391 430218 315711 430227
rect 37396 411903 165398 427903
rect 145398 409147 165398 411903
rect 145398 401839 146500 409147
rect 164068 401839 165398 409147
rect 315391 404023 315407 430218
rect 315644 404023 315711 430218
rect 315391 404007 315711 404023
rect 145398 400903 165398 401839
rect 363221 388853 364263 390887
rect 333727 388772 364263 388853
rect 333727 387884 333824 388772
rect 336416 387884 364263 388772
rect 333727 387811 364263 387884
<< via4 >>
rect 146520 674731 164088 681965
rect 178294 673993 192634 681741
rect 510140 694218 525390 700140
rect 146784 556095 164076 567969
rect 329310 625656 329890 666846
rect 443952 669616 462134 679662
rect 472834 676484 491834 680688
rect 327010 615420 327590 625656
rect 472272 599798 489906 613524
rect 350660 455969 355612 460921
rect 380103 451299 385103 456299
rect 146500 401839 164068 409147
rect 315407 404023 315496 430218
rect 315496 404023 315644 430218
rect 335540 391085 335860 391213
rect 335540 391021 335668 391085
rect 335668 391021 335732 391085
rect 335732 391021 335860 391085
rect 335540 390893 335860 391021
rect 334540 390151 334860 390274
rect 334540 390077 334663 390151
rect 334663 390077 334737 390151
rect 334737 390077 334860 390151
rect 334540 389954 334860 390077
<< metal5 >>
rect 509482 700140 525794 700828
rect 199140 694994 200140 700140
rect 199140 693994 215608 694994
rect 217076 694329 313018 700140
rect 217076 694064 326008 694329
rect 214608 686056 215608 693994
rect 303443 685915 326008 694064
rect 145394 681965 165394 682901
rect 145394 674731 146520 681965
rect 164088 674731 165394 681965
rect 145394 672901 165394 674731
rect 177396 681741 193396 682901
rect 177396 673993 178294 681741
rect 192634 673993 193396 681741
rect 177396 672901 193396 673993
rect 37396 655903 301396 671903
rect 318008 668449 326008 685915
rect 329491 680766 333977 700140
rect 344882 694218 510140 700140
rect 525390 694218 525836 700140
rect 344882 694016 525836 694218
rect 329491 669335 333996 680766
rect 344882 679466 352882 694016
rect 422585 692424 428028 694016
rect 509588 693836 525836 694016
rect 419347 680730 454676 683321
rect 472300 680730 492300 680984
rect 419347 680128 462918 680730
rect 344618 671466 352882 679466
rect 318008 667405 326803 668449
rect 318008 667076 329224 667405
rect 318008 666846 330218 667076
rect 37396 427903 53396 655903
rect 54394 638901 284394 654901
rect 54394 444901 70394 638901
rect 71394 621901 267394 637901
rect 71394 461901 87394 621901
rect 88394 604901 250394 620901
rect 88394 478901 104394 604901
rect 105394 587901 233394 604017
rect 105394 495901 121394 587901
rect 122394 567969 165394 569901
rect 122394 556095 146784 567969
rect 164076 556095 165394 567969
rect 122394 553901 165394 556095
rect 122394 512901 138394 553901
rect 217394 512901 233394 587901
rect 122394 496901 233394 512901
rect 234394 495901 250394 604901
rect 105394 479901 250394 495901
rect 251394 478901 267394 621901
rect 88394 462901 267394 478901
rect 268394 461901 284394 638901
rect 71394 445901 284394 461901
rect 285394 444901 301394 655903
rect 318008 641449 329310 666846
rect 320810 625656 329310 641449
rect 329890 625656 330218 666846
rect 333349 625826 333996 669335
rect 344882 650788 352882 671466
rect 442918 679662 462918 680128
rect 442918 669616 443952 679662
rect 462134 669616 462918 679662
rect 442918 668730 462918 669616
rect 470918 680688 492300 680730
rect 470918 676484 472834 680688
rect 491834 676484 492300 680688
rect 470918 675984 492300 676484
rect 470918 665730 490918 675984
rect 470918 649730 567918 665730
rect 365918 632730 550918 648730
rect 320810 615420 327010 625656
rect 327590 625550 330218 625656
rect 327590 615420 327934 625550
rect 320810 614586 327934 615420
rect 320810 595474 325810 614586
rect 320810 590474 338214 595474
rect 333214 460945 338214 590474
rect 365918 483730 381918 632730
rect 382918 615730 533918 631730
rect 382918 500730 398918 615730
rect 399918 613524 490918 614730
rect 399918 599798 472272 613524
rect 489906 599798 490918 613524
rect 399918 598730 490918 599798
rect 399918 517730 415918 598730
rect 517918 517730 533918 615730
rect 399918 501730 533918 517730
rect 534918 500730 550918 632730
rect 382918 484730 550918 500730
rect 551918 483730 567918 649730
rect 365918 467730 567918 483730
rect 333214 460921 355636 460945
rect 333214 455969 350660 460921
rect 355612 455969 355636 460921
rect 333214 455945 355636 455969
rect 361201 458168 571624 459210
rect 333214 454104 338214 455945
rect 54394 428901 301394 444901
rect 315381 453776 338214 454104
rect 315381 453774 332876 453776
rect 315381 430218 315711 453774
rect 361201 448109 362243 458168
rect 380079 456299 385127 456323
rect 380079 451299 380103 456299
rect 385103 451299 385127 456299
rect 380079 451275 385127 451299
rect 380103 450246 385103 451275
rect 380103 445246 411181 450246
rect 37396 411903 165398 427903
rect 145398 409147 165398 411903
rect 145398 401839 146500 409147
rect 164068 401839 165398 409147
rect 315381 404023 315407 430218
rect 315644 404023 315711 430218
rect 315381 403997 315711 404023
rect 145398 400903 165398 401839
rect 35194 391213 338981 391482
rect 35194 391026 335540 391213
rect 335516 390893 335540 391026
rect 335860 391026 338981 391213
rect 335860 390893 335884 391026
rect 335516 390869 335884 390893
rect 339620 390402 340085 392808
rect 35194 390274 340085 390402
rect 35194 389954 334540 390274
rect 334860 389954 340085 390274
rect 35194 389937 340085 389954
rect 334516 389930 334884 389937
<< comment >>
rect 528592 704000 564228 704100
use LDO  LDO_0
timestamp 1667842615
transform -1 0 550078 0 -1 694876
box -8958 -8682 15320 8530
use decoupling_cell  decoupling_cell_0
timestamp 1667074381
transform 1 0 368582 0 1 242038
box 0 0 201600 203879
use mirrors  mirrors_0
timestamp 1667846787
transform 0 -1 358618 1 0 616664
box -18962 22 70826 31618
use pwm_lower  pwm_lower_0
timestamp 1667170575
transform 0 1 413660 -1 0 697163
box 4398 -2478 18637 19086
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_0
timestamp 1667857442
transform 1 0 335699 0 1 389400
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_1
timestamp 1667857442
transform 1 0 334699 0 1 389400
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_2
timestamp 1667857442
transform 1 0 468123 0 1 450054
box -423 -423 423 423
use sky130_fd_pr__diode_pd2nw_11v0_K4SERG  sky130_fd_pr__diode_pd2nw_11v0_K4SERG_3
timestamp 1667857442
transform 1 0 469123 0 1 450054
box -423 -423 423 423
use switched_cap  switched_cap_0
timestamp 1667842615
transform -1 0 358010 0 -1 391814
box -6253 -57972 42538 2189
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
