magic
tech sky130A
magscale 1 2
timestamp 1665559092
<< pwell >>
rect -328 -823 328 823
<< mvnmos >>
rect -100 365 100 565
rect -100 55 100 255
rect -100 -255 100 -55
rect -100 -565 100 -365
<< mvndiff >>
rect -158 553 -100 565
rect -158 377 -146 553
rect -112 377 -100 553
rect -158 365 -100 377
rect 100 553 158 565
rect 100 377 112 553
rect 146 377 158 553
rect 100 365 158 377
rect -158 243 -100 255
rect -158 67 -146 243
rect -112 67 -100 243
rect -158 55 -100 67
rect 100 243 158 255
rect 100 67 112 243
rect 146 67 158 243
rect 100 55 158 67
rect -158 -67 -100 -55
rect -158 -243 -146 -67
rect -112 -243 -100 -67
rect -158 -255 -100 -243
rect 100 -67 158 -55
rect 100 -243 112 -67
rect 146 -243 158 -67
rect 100 -255 158 -243
rect -158 -377 -100 -365
rect -158 -553 -146 -377
rect -112 -553 -100 -377
rect -158 -565 -100 -553
rect 100 -377 158 -365
rect 100 -553 112 -377
rect 146 -553 158 -377
rect 100 -565 158 -553
<< mvndiffc >>
rect -146 377 -112 553
rect 112 377 146 553
rect -146 67 -112 243
rect 112 67 146 243
rect -146 -243 -112 -67
rect 112 -243 146 -67
rect -146 -553 -112 -377
rect 112 -553 146 -377
<< mvpsubdiff >>
rect -292 775 292 787
rect -292 741 -184 775
rect 184 741 292 775
rect -292 729 292 741
rect -292 679 -234 729
rect -292 -679 -280 679
rect -246 -679 -234 679
rect 234 679 292 729
rect -292 -729 -234 -679
rect 234 -679 246 679
rect 280 -679 292 679
rect 234 -729 292 -679
rect -292 -741 292 -729
rect -292 -775 -184 -741
rect 184 -775 292 -741
rect -292 -787 292 -775
<< mvpsubdiffcont >>
rect -184 741 184 775
rect -280 -679 -246 679
rect 246 -679 280 679
rect -184 -775 184 -741
<< poly >>
rect -100 637 100 653
rect -100 603 -84 637
rect 84 603 100 637
rect -100 565 100 603
rect -100 327 100 365
rect -100 293 -84 327
rect 84 293 100 327
rect -100 255 100 293
rect -100 17 100 55
rect -100 -17 -84 17
rect 84 -17 100 17
rect -100 -55 100 -17
rect -100 -293 100 -255
rect -100 -327 -84 -293
rect 84 -327 100 -293
rect -100 -365 100 -327
rect -100 -603 100 -565
rect -100 -637 -84 -603
rect 84 -637 100 -603
rect -100 -653 100 -637
<< polycont >>
rect -84 603 84 637
rect -84 293 84 327
rect -84 -17 84 17
rect -84 -327 84 -293
rect -84 -637 84 -603
<< locali >>
rect -280 741 -184 775
rect 184 741 280 775
rect -280 679 -246 741
rect 246 679 280 741
rect -100 603 -84 637
rect 84 603 100 637
rect -146 553 -112 569
rect -146 361 -112 377
rect 112 553 146 569
rect 112 361 146 377
rect -100 293 -84 327
rect 84 293 100 327
rect -146 243 -112 259
rect -146 51 -112 67
rect 112 243 146 259
rect 112 51 146 67
rect -100 -17 -84 17
rect 84 -17 100 17
rect -146 -67 -112 -51
rect -146 -259 -112 -243
rect 112 -67 146 -51
rect 112 -259 146 -243
rect -100 -327 -84 -293
rect 84 -327 100 -293
rect -146 -377 -112 -361
rect -146 -569 -112 -553
rect 112 -377 146 -361
rect 112 -569 146 -553
rect -100 -637 -84 -603
rect 84 -637 100 -603
rect -280 -741 -246 -679
rect 246 -741 280 -679
rect -280 -775 -184 -741
rect 184 -775 280 -741
<< viali >>
rect -84 603 84 637
rect -146 377 -112 553
rect 112 377 146 553
rect -84 293 84 327
rect -146 67 -112 243
rect 112 67 146 243
rect -84 -17 84 17
rect -146 -243 -112 -67
rect 112 -243 146 -67
rect -84 -327 84 -293
rect -146 -553 -112 -377
rect 112 -553 146 -377
rect -84 -637 84 -603
<< metal1 >>
rect -96 637 96 643
rect -96 603 -84 637
rect 84 603 96 637
rect -96 597 96 603
rect -152 553 -106 565
rect -152 377 -146 553
rect -112 377 -106 553
rect -152 365 -106 377
rect 106 553 152 565
rect 106 377 112 553
rect 146 377 152 553
rect 106 365 152 377
rect -96 327 96 333
rect -96 293 -84 327
rect 84 293 96 327
rect -96 287 96 293
rect -152 243 -106 255
rect -152 67 -146 243
rect -112 67 -106 243
rect -152 55 -106 67
rect 106 243 152 255
rect 106 67 112 243
rect 146 67 152 243
rect 106 55 152 67
rect -96 17 96 23
rect -96 -17 -84 17
rect 84 -17 96 17
rect -96 -23 96 -17
rect -152 -67 -106 -55
rect -152 -243 -146 -67
rect -112 -243 -106 -67
rect -152 -255 -106 -243
rect 106 -67 152 -55
rect 106 -243 112 -67
rect 146 -243 152 -67
rect 106 -255 152 -243
rect -96 -293 96 -287
rect -96 -327 -84 -293
rect 84 -327 96 -293
rect -96 -333 96 -327
rect -152 -377 -106 -365
rect -152 -553 -146 -377
rect -112 -553 -106 -377
rect -152 -565 -106 -553
rect 106 -377 152 -365
rect 106 -553 112 -377
rect 146 -553 152 -377
rect 106 -565 152 -553
rect -96 -603 96 -597
rect -96 -637 -84 -603
rect 84 -637 96 -603
rect -96 -643 96 -637
<< properties >>
string FIXED_BBOX -263 -758 263 758
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 1 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
