magic
tech sky130A
magscale 1 2
timestamp 1666558548
<< viali >>
rect -3254 5176 -3216 5212
rect -2604 5176 -2566 5212
rect -1958 5174 -1920 5210
rect -1250 5174 -1212 5210
rect -508 5174 -470 5210
rect 360 5174 398 5210
rect 1288 5174 1326 5210
rect 1794 5176 1832 5212
rect 2404 5176 2442 5212
rect 2946 5176 2984 5212
rect 3618 5176 3656 5212
rect 5092 5176 5130 5212
rect 6004 5178 6042 5214
rect 6696 5176 6734 5212
rect 7642 5176 7680 5212
rect 8182 5176 8220 5212
rect 8508 5176 8546 5212
rect 9142 5172 9180 5208
rect 1918 3838 1956 3874
rect 2204 3840 2242 3876
rect 2706 3840 2744 3876
rect 2980 3838 3018 3874
rect 3696 3836 3734 3872
rect 4142 3836 4180 3872
rect 4474 3838 4512 3874
rect 602 3728 640 3764
rect 864 3728 902 3764
rect 1170 3728 1208 3764
rect 1912 3722 1950 3758
rect 2202 3722 2240 3758
rect 2698 3722 2736 3758
rect 2976 3722 3014 3758
rect 3692 3724 3730 3760
rect 4140 3722 4178 3758
rect 4474 3720 4512 3756
rect 5056 3718 5094 3754
rect 5464 3718 5502 3754
rect 6010 3718 6048 3754
<< metal1 >>
rect 9358 5292 9558 5362
rect -3268 5212 -3206 5224
rect -3268 5176 -3254 5212
rect -3216 5176 -3206 5212
rect -3268 5118 -3206 5176
rect -2616 5212 -2554 5224
rect -2616 5176 -2604 5212
rect -2566 5176 -2554 5212
rect -2616 5118 -2554 5176
rect -1972 5210 -1910 5222
rect -1972 5174 -1958 5210
rect -1920 5174 -1910 5210
rect -1972 5118 -1910 5174
rect -1262 5210 -1200 5222
rect -1262 5174 -1250 5210
rect -1212 5174 -1200 5210
rect -1262 5118 -1200 5174
rect -522 5210 -460 5222
rect -522 5174 -508 5210
rect -470 5174 -460 5210
rect -522 5118 -460 5174
rect 348 5210 410 5222
rect 348 5174 360 5210
rect 398 5174 410 5210
rect 348 5118 410 5174
rect 1274 5210 1336 5222
rect 1274 5174 1288 5210
rect 1326 5174 1336 5210
rect 1274 5118 1336 5174
rect 1782 5212 1844 5224
rect 1782 5176 1794 5212
rect 1832 5176 1844 5212
rect 1782 5118 1844 5176
rect 2392 5212 2454 5222
rect 2392 5176 2404 5212
rect 2442 5176 2454 5212
rect 2392 5118 2454 5176
rect 2934 5212 2996 5224
rect 2934 5176 2946 5212
rect 2984 5176 2996 5212
rect 2934 5118 2996 5176
rect 3606 5212 3668 5224
rect 3606 5176 3618 5212
rect 3656 5176 3668 5212
rect 3606 5118 3668 5176
rect 5078 5212 5148 5226
rect 5078 5176 5092 5212
rect 5130 5176 5148 5212
rect 5078 5118 5148 5176
rect 5988 5214 6056 5226
rect 5988 5178 6004 5214
rect 6042 5178 6056 5214
rect 5988 5118 6056 5178
rect 6682 5212 6752 5224
rect 6682 5176 6696 5212
rect 6734 5176 6752 5212
rect 6682 5118 6752 5176
rect 7626 5212 7696 5226
rect 7626 5176 7642 5212
rect 7680 5176 7696 5212
rect 7626 5118 7696 5176
rect 8168 5212 8238 5224
rect 8168 5176 8182 5212
rect 8220 5176 8238 5212
rect 8168 5118 8238 5176
rect 8496 5212 8558 5222
rect 8496 5176 8508 5212
rect 8546 5176 8558 5212
rect 8496 5118 8558 5176
rect 9130 5208 9200 5224
rect 9130 5172 9142 5208
rect 9180 5172 9200 5208
rect 9130 5118 9200 5172
rect 9424 5118 9486 5292
rect -3536 5068 9486 5118
rect -3536 5066 -3390 5068
rect -3538 4904 4664 4954
rect 4778 4906 9736 4956
rect -3838 4806 -3774 4812
rect -3838 4754 -3832 4806
rect -3780 4756 4436 4806
rect 4614 4792 4664 4904
rect 7652 4798 7702 4906
rect 8130 4798 8180 4906
rect 8682 4798 8732 4906
rect 9192 4798 9242 4906
rect -3780 4754 -3774 4756
rect -3838 4748 -3774 4754
rect -3580 4644 -3530 4756
rect 4614 4742 6954 4792
rect 7214 4750 9506 4798
rect -3580 4596 -3032 4644
rect -3300 4560 -3032 4596
rect -3272 4556 -3068 4560
rect -3272 4440 -3260 4556
rect -3080 4440 -3068 4556
rect 1268 4540 1332 4544
rect 1268 4488 1274 4540
rect 1326 4534 1332 4540
rect 4614 4534 4664 4742
rect 1326 4488 4664 4534
rect 6610 4550 6674 4556
rect 7214 4550 7264 4750
rect 6610 4548 7264 4550
rect 6610 4496 6618 4548
rect 6670 4500 7264 4548
rect 6670 4496 6674 4500
rect 7214 4498 7264 4500
rect 6610 4488 6674 4496
rect 1268 4484 4664 4488
rect 1268 4476 1332 4484
rect -3272 4428 -3068 4440
rect 6372 4304 6434 4312
rect 1768 4302 6434 4304
rect 1768 4254 6378 4302
rect 6372 4250 6378 4254
rect 6430 4250 6434 4302
rect 6372 4244 6434 4250
rect 5178 4154 5244 4162
rect 1518 4146 1584 4154
rect 1518 4094 1524 4146
rect 1576 4144 1584 4146
rect 5178 4144 5184 4154
rect 1576 4094 3250 4144
rect 3530 4102 5184 4144
rect 5236 4102 5244 4154
rect 3530 4094 5244 4102
rect 1518 4086 1584 4094
rect 1270 3992 1334 4000
rect 1270 3940 1276 3992
rect 1328 3990 1334 3992
rect 6612 3996 6676 4002
rect 6612 3990 6618 3996
rect 1328 3940 3284 3990
rect 3440 3944 6618 3990
rect 6670 3944 6676 3996
rect 3440 3940 6676 3944
rect 1270 3932 1334 3940
rect 6612 3934 6676 3940
rect 1890 3874 1974 3884
rect 1890 3838 1918 3874
rect 1956 3838 1974 3874
rect 586 3764 658 3778
rect 586 3728 602 3764
rect 640 3728 658 3764
rect 586 3664 658 3728
rect 850 3764 922 3778
rect 850 3728 864 3764
rect 902 3728 922 3764
rect 850 3664 922 3728
rect 1150 3764 1222 3778
rect 1150 3728 1170 3764
rect 1208 3728 1222 3764
rect 1150 3664 1222 3728
rect 1890 3758 1974 3838
rect 1890 3722 1912 3758
rect 1950 3722 1974 3758
rect 1890 3664 1974 3722
rect 2182 3876 2266 3886
rect 2182 3840 2204 3876
rect 2242 3840 2266 3876
rect 2182 3758 2266 3840
rect 2182 3722 2202 3758
rect 2240 3722 2266 3758
rect 2182 3664 2266 3722
rect 2686 3876 2770 3886
rect 2686 3840 2706 3876
rect 2744 3840 2770 3876
rect 2686 3758 2770 3840
rect 2686 3722 2698 3758
rect 2736 3722 2770 3758
rect 2686 3664 2770 3722
rect 2954 3874 3036 3884
rect 2954 3838 2980 3874
rect 3018 3838 3036 3874
rect 2954 3758 3036 3838
rect 2954 3722 2976 3758
rect 3014 3722 3036 3758
rect 2954 3664 3036 3722
rect 3678 3872 3754 3884
rect 3678 3836 3696 3872
rect 3734 3836 3754 3872
rect 3678 3760 3754 3836
rect 3678 3724 3692 3760
rect 3730 3724 3754 3760
rect 3678 3664 3754 3724
rect 4120 3872 4196 3884
rect 4120 3836 4142 3872
rect 4180 3836 4196 3872
rect 4120 3758 4196 3836
rect 4120 3722 4140 3758
rect 4178 3722 4196 3758
rect 4120 3664 4196 3722
rect 4456 3874 4532 3882
rect 4456 3838 4474 3874
rect 4512 3838 4532 3874
rect 4456 3756 4532 3838
rect 4456 3720 4474 3756
rect 4512 3720 4532 3756
rect 4456 3664 4532 3720
rect 5046 3754 5100 3766
rect 5046 3718 5056 3754
rect 5094 3718 5100 3754
rect 5046 3664 5100 3718
rect 5456 3754 5510 3766
rect 5456 3718 5464 3754
rect 5502 3718 5510 3754
rect 5456 3664 5510 3718
rect 6000 3754 6054 3766
rect 6000 3718 6010 3754
rect 6048 3718 6054 3754
rect 6000 3664 6054 3718
rect 6536 3664 6606 3732
rect 312 3614 6606 3664
rect 6536 3532 6606 3614
rect 288 3448 6188 3498
rect -3838 3360 -3774 3366
rect -3838 3308 -3832 3360
rect -3780 3356 -3774 3360
rect -3780 3308 1346 3356
rect 2338 3348 2390 3448
rect 2648 3348 2700 3448
rect -3838 3304 1346 3308
rect -3838 3298 -3774 3304
rect 1766 3298 4566 3348
rect 6372 3340 6434 3348
rect 6372 3338 6378 3340
rect 3230 3148 3280 3298
rect 4908 3288 6378 3338
rect 6430 3288 6434 3340
rect 6372 3282 6434 3288
<< via1 >>
rect -3832 4754 -3780 4806
rect -3260 4440 -3080 4556
rect 1274 4488 1326 4540
rect 6618 4496 6670 4548
rect 6378 4250 6430 4302
rect 1524 4094 1576 4146
rect 5184 4102 5236 4154
rect 1276 3940 1328 3992
rect 6618 3944 6670 3996
rect -3832 3308 -3780 3360
rect 6378 3288 6430 3340
<< metal2 >>
rect 1452 6088 1652 6158
rect 5112 6096 5312 6166
rect -3838 4806 -3774 4812
rect -3838 4754 -3832 4806
rect -3780 4754 -3774 4806
rect -3838 4748 -3774 4754
rect -3832 4398 -3780 4748
rect -3286 4562 -3068 4574
rect -3286 4432 -3272 4562
rect -3084 4556 -3068 4562
rect -3080 4440 -3068 4556
rect 1268 4540 1332 4544
rect 1268 4488 1274 4540
rect 1326 4488 1332 4540
rect 1268 4476 1332 4488
rect -3084 4432 -3068 4440
rect -3286 4420 -3068 4432
rect -4388 4348 -3780 4398
rect 1276 4378 1326 4476
rect -3832 3366 -3780 4348
rect -284 4338 1326 4378
rect -284 4328 -256 4338
rect -268 4266 -256 4328
rect -186 4328 1326 4338
rect -186 4266 -170 4328
rect -268 4254 -170 4266
rect 1276 4000 1326 4328
rect 1524 4154 1574 6088
rect 5184 4162 5234 6096
rect 6610 4548 6674 4556
rect 6610 4496 6618 4548
rect 6670 4496 6674 4548
rect 6610 4488 6674 4496
rect 6372 4302 6434 4312
rect 6372 4250 6378 4302
rect 6430 4250 6434 4302
rect 6372 4244 6434 4250
rect 5178 4154 5244 4162
rect 1518 4146 1584 4154
rect 1518 4094 1524 4146
rect 1576 4094 1584 4146
rect 5178 4102 5184 4154
rect 5236 4102 5244 4154
rect 5178 4094 5244 4102
rect 1518 4086 1584 4094
rect 1270 3992 1334 4000
rect 1270 3940 1276 3992
rect 1328 3940 1334 3992
rect 1270 3932 1334 3940
rect -3838 3360 -3774 3366
rect -3838 3308 -3832 3360
rect -3780 3308 -3774 3360
rect 6378 3348 6428 4244
rect 6618 4002 6668 4488
rect 6612 3996 6676 4002
rect 6612 3944 6618 3996
rect 6670 3944 6676 3996
rect 6612 3934 6676 3944
rect -3838 3298 -3774 3308
rect 6372 3340 6434 3348
rect 6372 3288 6378 3340
rect 6430 3288 6434 3340
rect 6372 3282 6434 3288
<< via2 >>
rect -3272 4556 -3084 4562
rect -3272 4440 -3260 4556
rect -3260 4440 -3084 4556
rect -3272 4432 -3084 4440
rect -256 4266 -186 4338
<< metal3 >>
rect -3310 4576 -3036 4584
rect -3310 4418 -3292 4576
rect -3056 4418 -3036 4576
rect -3310 4408 -3036 4418
rect -272 4346 -170 4354
rect -272 4258 -264 4346
rect -178 4258 -170 4346
rect -272 4250 -170 4258
<< via3 >>
rect -3292 4562 -3056 4576
rect -3292 4432 -3272 4562
rect -3272 4432 -3084 4562
rect -3084 4432 -3056 4562
rect -3292 4418 -3056 4432
rect -264 4338 -178 4346
rect -264 4266 -256 4338
rect -256 4266 -186 4338
rect -186 4266 -178 4338
rect -264 4258 -178 4266
<< metal4 >>
rect -284 4346 -154 4378
rect -284 4258 -264 4346
rect -178 4258 -154 4346
rect -284 4224 -154 4258
<< via4 >>
rect -3372 4576 -2972 4612
rect -3372 4418 -3292 4576
rect -3292 4418 -3056 4576
rect -3056 4418 -2972 4576
rect -3372 4370 -2972 4418
<< metal5 >>
rect -3396 4612 -2942 4644
rect -3396 4370 -3372 4612
rect -2972 4370 -2942 4612
rect -3396 3930 -2942 4370
use sky130_fd_pr__cap_mim_m3_2_GH5TRZ  sky130_fd_pr__cap_mim_m3_2_GH5TRZ_0
timestamp 1665683293
transform 1 0 -1922 0 1 2770
box -1766 -1516 1788 1516
use sky130_fd_pr__nfet_g5v0d10v5_8PFU4A  sky130_fd_pr__nfet_g5v0d10v5_8PFU4A_0
timestamp 1665559092
transform 0 1 888 -1 0 3482
box -328 -668 328 668
use sky130_fd_pr__nfet_g5v0d10v5_FEGU4A  sky130_fd_pr__nfet_g5v0d10v5_FEGU4A_0
timestamp 1665559092
transform 0 1 5553 -1 0 3472
box -328 -823 328 823
use sky130_fd_pr__nfet_g5v0d10v5_FEGU4A  sky130_fd_pr__nfet_g5v0d10v5_FEGU4A_1
timestamp 1665559092
transform 0 1 2545 -1 0 4118
box -328 -823 328 823
use sky130_fd_pr__nfet_g5v0d10v5_FEGU4A  sky130_fd_pr__nfet_g5v0d10v5_FEGU4A_2
timestamp 1665559092
transform 0 1 4175 -1 0 4116
box -328 -823 328 823
use sky130_fd_pr__nfet_g5v0d10v5_NQKU4A  sky130_fd_pr__nfet_g5v0d10v5_NQKU4A_0
timestamp 1665559092
transform 0 1 3140 -1 0 3476
box -328 -1598 328 1598
use sky130_fd_pr__pfet_g5v0d10v5_2JCT5W  sky130_fd_pr__pfet_g5v0d10v5_2JCT5W_0
timestamp 1665560597
transform 0 -1 477 1 0 4930
box -358 -4193 358 4193
use sky130_fd_pr__pfet_g5v0d10v5_QS9L5N  sky130_fd_pr__pfet_g5v0d10v5_QS9L5N_0
timestamp 1665560017
transform 0 1 8449 -1 0 4930
box -358 -1289 358 1289
use sky130_fd_pr__pfet_g5v0d10v5_QS9L5N  sky130_fd_pr__pfet_g5v0d10v5_QS9L5N_1
timestamp 1665560017
transform 0 1 5893 -1 0 4930
box -358 -1289 358 1289
<< labels >>
rlabel metal1 6552 3558 6592 3716 1 Vminus
rlabel metal1 9376 5308 9532 5348 1 Vplus
rlabel metal2 5128 6110 5284 6150 1 Vin1
rlabel metal2 1476 6102 1632 6142 1 Vin2
rlabel metal2 -4378 4358 -4330 4384 1 Out
<< end >>
