magic
tech sky130A
magscale 1 2
timestamp 1665943203
<< locali >>
rect -268 1860 634 1894
rect -268 1700 -234 1860
rect -268 1130 -120 1700
rect -268 986 -234 1130
rect 600 986 634 1860
rect 1314 1860 2216 1894
rect 1314 1700 1348 1860
rect 1314 1130 1462 1700
rect 2182 1130 2216 1860
rect 1314 986 1348 1130
rect 2182 1096 3760 1130
rect 5574 1096 5670 1130
rect 2182 986 2216 1096
rect -268 952 2216 986
rect -20 832 76 866
rect 1134 832 1422 866
rect 2482 832 2578 866
rect -20 498 14 832
rect -424 464 -328 498
rect -190 464 14 498
rect -424 402 -390 464
rect -424 -238 -390 64
rect -128 402 14 464
rect -94 52 14 402
rect -128 -120 14 52
rect 1196 -120 1362 832
rect 2542 770 2578 832
rect 2542 -58 2544 770
rect 2578 114 2760 148
rect 3310 114 3406 148
rect 2578 -22 2698 114
rect 3372 52 3406 114
rect 2578 -58 2812 -22
rect 2542 -120 2812 -58
rect -128 -154 1482 -120
rect 2482 -154 2812 -120
rect -128 -220 1574 -154
rect -94 -226 1574 -220
rect -94 -228 888 -226
rect -424 -742 -390 -680
rect -94 -262 76 -228
rect 626 -262 888 -228
rect 1442 -262 1574 -226
rect -94 -324 14 -262
rect -94 -362 -20 -324
rect -94 -364 14 -362
rect -128 -642 14 -364
rect 688 -398 829 -262
rect 1503 -398 1574 -262
rect 574 -606 829 -398
rect 1388 -606 1574 -398
rect -128 -680 -20 -642
rect -128 -742 14 -680
rect 318 -684 382 -640
rect 688 -742 829 -606
rect 1503 -708 1574 -606
rect 2664 -408 2812 -154
rect 2698 -600 2812 -408
rect 2664 -606 2812 -600
rect 2664 -708 2698 -606
rect 1503 -742 2698 -708
rect 3488 -676 3522 1096
rect 5636 1034 5670 1096
rect 5636 -642 5670 -580
rect 3536 -676 3584 -642
rect 5574 -676 5670 -642
rect 3372 -742 3406 -680
rect -424 -776 -328 -742
rect -190 -776 76 -742
rect 596 -776 994 -742
rect 1352 -776 2882 -742
rect 3196 -776 3406 -742
<< viali >>
rect 3760 1096 5574 1130
rect 76 832 1134 866
rect 1422 832 2482 866
rect -328 464 -190 498
rect -424 64 -390 402
rect -128 52 -94 402
rect 2544 -58 2578 770
rect 2760 114 3310 148
rect 1482 -154 2482 -120
rect -424 -680 -390 -238
rect -128 -364 -94 -228
rect 76 -262 626 -228
rect 888 -262 1442 -226
rect -20 -362 14 -324
rect -20 -680 14 -642
rect 2664 -600 2698 -408
rect 3372 -680 3406 52
rect 5636 -580 5670 1034
rect 3584 -676 5574 -642
rect -328 -776 -190 -742
rect 76 -776 596 -742
rect 994 -776 1352 -742
rect 2882 -776 3196 -742
<< metal1 >>
rect 18 1848 30 1906
rect 328 1848 340 1906
rect 1594 1848 1606 1906
rect 1904 1848 1916 1906
rect -108 1752 2056 1808
rect 2912 1780 3396 1790
rect -32 1706 14 1752
rect 224 1706 270 1752
rect 480 1706 526 1752
rect -178 1700 -114 1706
rect -178 1146 -172 1700
rect -120 1146 -114 1700
rect -178 1140 -114 1146
rect -42 1700 24 1706
rect -42 1146 -36 1700
rect 18 1146 24 1700
rect -42 1140 24 1146
rect 90 1700 148 1706
rect 90 1146 92 1700
rect 146 1146 148 1700
rect 90 1140 148 1146
rect 214 1700 280 1706
rect 214 1146 220 1700
rect 274 1146 280 1700
rect 214 1140 280 1146
rect 346 1700 404 1706
rect 346 1146 348 1700
rect 402 1146 404 1700
rect 346 1140 404 1146
rect 470 1700 536 1706
rect 470 1146 476 1700
rect 530 1146 536 1700
rect 470 1140 536 1146
rect 1404 1700 1468 1706
rect 1404 1146 1410 1700
rect 1462 1146 1468 1700
rect 1404 1140 1468 1146
rect 1540 1700 1606 1706
rect 1540 1146 1546 1700
rect 1600 1146 1606 1700
rect 1540 1140 1606 1146
rect 1668 1700 1734 1706
rect 1668 1146 1674 1700
rect 1728 1146 1734 1700
rect 1668 1140 1734 1146
rect 1796 1700 1862 1706
rect 1796 1146 1802 1700
rect 1856 1146 1862 1700
rect 1796 1140 1862 1146
rect 1924 1700 1990 1706
rect 1924 1146 1930 1700
rect 1984 1146 1990 1700
rect 1924 1140 1990 1146
rect 2052 1700 2118 1706
rect 2052 1146 2058 1700
rect 2112 1146 2118 1700
rect 2052 1140 2118 1146
rect 2912 1494 2922 1780
rect 3386 1494 3396 1780
rect -32 1094 14 1140
rect 224 1094 270 1140
rect 480 1094 526 1140
rect -108 1038 2056 1094
rect 2912 1044 3396 1494
rect 3684 1140 4830 1142
rect 3684 1086 3696 1140
rect 5532 1130 5682 1142
rect 5574 1096 5682 1130
rect 5532 1086 5682 1096
rect 2768 1004 5510 1044
rect 2768 918 2776 1004
rect 2876 988 5510 1004
rect 5626 1034 5682 1086
rect 2876 918 3534 988
rect 2768 912 3534 918
rect -170 866 2598 886
rect -170 832 76 866
rect 1134 832 1422 866
rect 2482 832 2598 866
rect -170 820 2598 832
rect -170 506 -104 820
rect 2522 770 2598 820
rect 2 688 1130 744
rect 1282 688 2396 744
rect -432 498 -82 506
rect -432 464 -328 498
rect -190 464 -82 498
rect -432 456 -82 464
rect -432 402 -382 456
rect -432 64 -424 402
rect -390 64 -382 402
rect -140 402 -82 456
rect -432 52 -382 64
rect -294 54 -286 368
rect -234 54 -224 368
rect -140 52 -128 402
rect -94 52 -82 402
rect -140 40 -82 52
rect 2 24 52 688
rect 266 650 312 656
rect 424 650 470 656
rect 582 650 628 656
rect 740 650 786 656
rect 898 650 944 656
rect 1056 650 1102 656
rect 98 644 164 650
rect 98 68 104 644
rect 158 68 164 644
rect 98 62 164 68
rect 256 644 322 650
rect 256 68 262 644
rect 316 68 322 644
rect 256 62 322 68
rect 414 644 480 650
rect 414 68 420 644
rect 474 68 480 644
rect 414 62 480 68
rect 572 644 638 650
rect 572 68 578 644
rect 632 68 638 644
rect 572 62 638 68
rect 730 644 796 650
rect 730 68 736 644
rect 790 68 796 644
rect 730 62 796 68
rect 888 644 954 650
rect 888 68 894 644
rect 948 68 954 644
rect 888 62 954 68
rect 1046 644 1112 650
rect 1046 68 1052 644
rect 1106 68 1112 644
rect 1046 62 1112 68
rect 266 56 312 62
rect 424 56 470 62
rect 582 56 628 62
rect 740 56 786 62
rect 898 56 944 62
rect 1056 56 1102 62
rect 1282 24 1374 688
rect 1444 644 1510 650
rect 1444 68 1450 644
rect 1504 68 1510 644
rect 1444 62 1510 68
rect 1602 644 1668 650
rect 1602 68 1608 644
rect 1662 68 1668 644
rect 1602 62 1668 68
rect 1760 644 1826 650
rect 1760 68 1766 644
rect 1820 68 1826 644
rect 1760 62 1826 68
rect 1918 644 1984 650
rect 1918 68 1924 644
rect 1978 68 1984 644
rect 1918 62 1984 68
rect 2076 644 2142 650
rect 2076 68 2082 644
rect 2136 68 2142 644
rect 2076 62 2142 68
rect 2234 644 2300 650
rect 2234 68 2240 644
rect 2294 68 2300 644
rect 2234 62 2300 68
rect 2392 644 2458 650
rect 2392 68 2398 644
rect 2452 68 2458 644
rect 2392 62 2458 68
rect 2 22 1050 24
rect -460 14 -388 22
rect -460 -62 -454 14
rect -394 -62 -388 14
rect -460 -68 -388 -62
rect -32 14 1050 22
rect -32 -62 -26 14
rect 46 -32 1050 14
rect 1282 -32 2396 24
rect 46 -62 52 -32
rect -32 -68 52 -62
rect 1282 -96 1374 -32
rect -460 -188 1374 -96
rect 2522 -58 2544 770
rect 2578 156 2598 770
rect 2578 148 3414 156
rect 2578 114 2760 148
rect 3310 114 3414 148
rect 2578 106 3414 114
rect 2578 -58 2598 106
rect 2522 -98 2598 -58
rect 1464 -120 2598 -98
rect 1464 -154 1482 -120
rect 2482 -154 2598 -120
rect 1464 -174 2598 -154
rect 2656 6 3164 62
rect 3364 52 3414 106
rect -140 -220 -82 -216
rect 1464 -220 1536 -174
rect -140 -226 650 -220
rect 880 -226 1536 -220
rect -438 -238 -374 -226
rect -438 -680 -424 -238
rect -390 -680 -374 -238
rect -140 -228 888 -226
rect -140 -364 -128 -228
rect -94 -262 76 -228
rect 626 -262 888 -228
rect 1442 -262 1536 -226
rect -94 -270 650 -262
rect 880 -270 1472 -262
rect -94 -364 -82 -270
rect -140 -374 -82 -364
rect -32 -324 34 -270
rect 2656 -314 2712 6
rect -32 -362 -20 -324
rect 14 -362 34 -324
rect -32 -374 34 -362
rect 82 -370 2712 -314
rect 2760 -38 2824 -32
rect 82 -402 134 -370
rect -294 -602 134 -402
rect 174 -414 240 -408
rect 174 -590 180 -414
rect 234 -590 240 -414
rect 174 -596 240 -590
rect -438 -726 -374 -680
rect -28 -642 22 -630
rect -28 -680 -20 -642
rect 14 -680 22 -642
rect -28 -726 22 -680
rect 82 -634 134 -602
rect 280 -634 326 -370
rect 366 -414 432 -408
rect 366 -590 372 -414
rect 426 -590 432 -414
rect 366 -596 432 -590
rect 472 -634 518 -370
rect 558 -414 624 -408
rect 558 -590 564 -414
rect 618 -590 624 -414
rect 558 -596 624 -590
rect 734 -634 782 -370
rect 892 -414 956 -408
rect 892 -590 898 -414
rect 950 -590 956 -414
rect 892 -596 956 -590
rect 988 -414 1054 -408
rect 988 -590 994 -414
rect 1048 -590 1054 -414
rect 988 -596 1054 -590
rect 1086 -414 1150 -408
rect 1086 -590 1092 -414
rect 1144 -590 1150 -414
rect 1086 -596 1150 -590
rect 1182 -414 1248 -408
rect 1182 -590 1188 -414
rect 1240 -590 1248 -414
rect 1182 -596 1248 -590
rect 1278 -414 1342 -408
rect 1278 -590 1284 -414
rect 1336 -590 1342 -414
rect 1278 -596 1342 -590
rect 1374 -414 1438 -408
rect 1374 -590 1380 -414
rect 1432 -590 1438 -414
rect 1374 -596 1438 -590
rect 1548 -634 1604 -370
rect 2760 -402 2766 -38
rect 2652 -408 2766 -402
rect 2652 -600 2664 -408
rect 2698 -590 2766 -408
rect 2818 -590 2824 -38
rect 2698 -600 2824 -590
rect 2860 -38 2924 -32
rect 2860 -590 2866 -38
rect 2918 -590 2924 -38
rect 2860 -596 2924 -590
rect 2956 -38 3020 -32
rect 2956 -590 2962 -38
rect 3014 -590 3020 -38
rect 2956 -596 3020 -590
rect 3052 -38 3116 -32
rect 3052 -590 3058 -38
rect 3110 -590 3116 -38
rect 3052 -596 3116 -590
rect 3148 -38 3212 -32
rect 3148 -590 3154 -38
rect 3206 -590 3212 -38
rect 3148 -596 3212 -590
rect 3244 -38 3308 -32
rect 3244 -590 3250 -38
rect 3302 -590 3308 -38
rect 3244 -596 3308 -590
rect 2652 -606 2824 -600
rect 82 -690 3260 -634
rect 3364 -680 3372 52
rect 3406 -680 3414 52
rect 3478 -534 3534 912
rect 3584 936 3648 942
rect 3584 -482 3590 936
rect 3642 -482 3648 936
rect 3714 936 3778 942
rect 3714 -482 3720 936
rect 3772 -482 3778 936
rect 3844 936 3908 942
rect 3844 -482 3850 936
rect 3902 -482 3908 936
rect 3970 936 4034 942
rect 3970 -482 3976 936
rect 4028 -482 4034 936
rect 4100 936 4164 942
rect 4100 -482 4106 936
rect 4158 -482 4164 936
rect 4226 936 4290 942
rect 4226 -482 4232 936
rect 4284 -482 4290 936
rect 4356 936 4420 942
rect 4356 -482 4362 936
rect 4414 -482 4420 936
rect 4482 936 4546 942
rect 4482 -482 4488 936
rect 4540 -482 4546 936
rect 4612 936 4676 942
rect 4612 -482 4618 936
rect 4670 -482 4676 936
rect 4738 936 4802 942
rect 4738 -482 4744 936
rect 4796 -482 4802 936
rect 4868 936 4932 942
rect 4868 -482 4874 936
rect 4926 -482 4932 936
rect 4994 936 5058 942
rect 4994 -482 5000 936
rect 5052 -482 5058 936
rect 5124 936 5188 942
rect 5124 -482 5130 936
rect 5182 -482 5188 936
rect 5250 936 5314 942
rect 5250 -482 5256 936
rect 5308 -482 5314 936
rect 5380 936 5444 942
rect 5380 -482 5386 936
rect 5438 -482 5444 936
rect 5506 936 5570 942
rect 5506 -482 5512 936
rect 5564 -482 5570 936
rect 3478 -590 5510 -534
rect 5626 -580 5636 1034
rect 5670 -580 5682 1034
rect 5626 -632 5682 -580
rect -438 -732 604 -726
rect -438 -742 240 -732
rect -438 -776 -328 -742
rect -190 -776 76 -742
rect -438 -784 240 -776
rect 596 -784 604 -732
rect -438 -790 604 -784
rect 988 -732 1358 -726
rect 3364 -728 3414 -680
rect 3536 -642 5682 -632
rect 3536 -676 3584 -642
rect 5574 -676 5682 -642
rect 3536 -688 5682 -676
rect 988 -784 994 -732
rect 1352 -784 1358 -732
rect 988 -790 1358 -784
rect 2812 -734 3414 -728
rect 2812 -788 2818 -734
rect 3250 -788 3414 -734
rect 2812 -794 3414 -788
<< via1 >>
rect 30 1848 328 1906
rect 1606 1848 1904 1906
rect -172 1146 -120 1700
rect -36 1146 18 1700
rect 92 1146 146 1700
rect 220 1146 274 1700
rect 348 1146 402 1700
rect 476 1146 530 1700
rect 1410 1146 1462 1700
rect 1546 1146 1600 1700
rect 1674 1146 1728 1700
rect 1802 1146 1856 1700
rect 1930 1146 1984 1700
rect 2058 1146 2112 1700
rect 2922 1494 3386 1780
rect 4830 1140 5532 1142
rect 3696 1130 5532 1140
rect 3696 1096 3760 1130
rect 3760 1096 5532 1130
rect 3696 1086 5532 1096
rect 2776 918 2876 1004
rect -286 54 -234 368
rect 104 68 158 644
rect 262 68 316 644
rect 420 68 474 644
rect 578 68 632 644
rect 736 68 790 644
rect 894 68 948 644
rect 1052 68 1106 644
rect 1450 68 1504 644
rect 1608 68 1662 644
rect 1766 68 1820 644
rect 1924 68 1978 644
rect 2082 68 2136 644
rect 2240 68 2294 644
rect 2398 68 2452 644
rect -454 -62 -394 14
rect -26 -62 46 14
rect 180 -590 234 -414
rect 372 -590 426 -414
rect 564 -590 618 -414
rect 898 -590 950 -414
rect 994 -590 1048 -414
rect 1092 -590 1144 -414
rect 1188 -590 1240 -414
rect 1284 -590 1336 -414
rect 1380 -590 1432 -414
rect 2766 -590 2818 -38
rect 2866 -590 2918 -38
rect 2962 -590 3014 -38
rect 3058 -590 3110 -38
rect 3154 -590 3206 -38
rect 3250 -590 3302 -38
rect 3590 -482 3642 936
rect 3720 -482 3772 936
rect 3850 -482 3902 936
rect 3976 -482 4028 936
rect 4106 -482 4158 936
rect 4232 -482 4284 936
rect 4362 -482 4414 936
rect 4488 -482 4540 936
rect 4618 -482 4670 936
rect 4744 -482 4796 936
rect 4874 -482 4926 936
rect 5000 -482 5052 936
rect 5130 -482 5182 936
rect 5256 -482 5308 936
rect 5386 -482 5438 936
rect 5512 -482 5564 936
rect 240 -742 596 -732
rect 240 -776 596 -742
rect 240 -784 596 -776
rect 994 -742 1352 -732
rect 994 -776 1352 -742
rect 994 -784 1352 -776
rect 2818 -742 3250 -734
rect 2818 -776 2882 -742
rect 2882 -776 3196 -742
rect 3196 -776 3250 -742
rect 2818 -788 3250 -776
<< metal2 >>
rect -178 1906 2252 1930
rect -178 1848 30 1906
rect 328 1848 1606 1906
rect 1904 1848 2252 1906
rect -178 1838 2252 1848
rect -178 1700 -114 1838
rect -178 1146 -172 1700
rect -120 1146 -114 1700
rect -178 828 -114 1146
rect -42 1700 24 1706
rect -42 1146 -36 1700
rect 18 1146 24 1700
rect -42 1008 24 1146
rect 90 1700 148 1838
rect 90 1146 92 1700
rect 146 1146 148 1700
rect 90 1140 148 1146
rect 214 1700 280 1706
rect 214 1146 220 1700
rect 274 1146 280 1700
rect 214 1008 280 1146
rect 346 1700 404 1838
rect 346 1146 348 1700
rect 402 1146 404 1700
rect 346 1140 404 1146
rect 470 1700 536 1706
rect 470 1146 476 1700
rect 530 1146 536 1700
rect 470 1008 536 1146
rect 1404 1700 1468 1838
rect 1404 1146 1410 1700
rect 1462 1146 1468 1700
rect 1404 1140 1468 1146
rect 1540 1700 1606 1706
rect 1540 1146 1546 1700
rect 1600 1146 1606 1700
rect 1540 1008 1606 1146
rect 1672 1700 1730 1838
rect 1672 1146 1674 1700
rect 1728 1146 1730 1700
rect 1672 1140 1730 1146
rect 1796 1700 1862 1706
rect 1796 1146 1802 1700
rect 1856 1146 1862 1700
rect 1796 1008 1862 1146
rect 1928 1700 1986 1838
rect 1928 1146 1930 1700
rect 1984 1146 1986 1700
rect 1928 1140 1986 1146
rect 2052 1700 2118 1706
rect 2052 1146 2058 1700
rect 2112 1146 2118 1700
rect 2052 1008 2118 1146
rect 2160 1244 2252 1838
rect 2912 1780 3396 1790
rect 2912 1494 2922 1780
rect 3386 1494 3396 1780
rect 2912 1484 3396 1494
rect 4036 1244 4636 1814
rect 2160 1142 5570 1244
rect 2160 1140 4830 1142
rect 2160 1086 3696 1140
rect 5532 1086 5570 1142
rect 2160 1068 5570 1086
rect -42 916 1112 1008
rect -292 764 -114 828
rect -292 368 -228 764
rect -292 54 -286 368
rect -234 54 -228 368
rect 98 644 164 916
rect 98 68 104 644
rect 158 68 164 644
rect 98 62 164 68
rect 256 644 322 656
rect 256 68 262 644
rect 316 68 322 644
rect -292 48 -228 54
rect -460 14 52 20
rect -460 -62 -454 14
rect -394 -62 -26 14
rect 46 -62 52 14
rect -460 -68 52 -62
rect 256 -44 322 68
rect 414 644 480 916
rect 414 68 420 644
rect 474 68 480 644
rect 414 62 480 68
rect 572 644 638 656
rect 572 68 578 644
rect 632 68 638 644
rect 572 -44 638 68
rect 730 644 796 916
rect 730 68 736 644
rect 790 68 796 644
rect 730 62 796 68
rect 888 644 954 656
rect 888 68 894 644
rect 948 68 954 644
rect 888 -44 954 68
rect 1046 644 1112 916
rect 1046 68 1052 644
rect 1106 68 1112 644
rect 1046 62 1112 68
rect 1444 1004 2882 1008
rect 1444 918 2776 1004
rect 2876 918 2882 1004
rect 1444 916 2882 918
rect 3584 936 3648 942
rect 1444 644 1510 916
rect 1444 68 1450 644
rect 1504 68 1510 644
rect 1444 62 1510 68
rect 1602 644 1668 650
rect 1602 68 1608 644
rect 1662 68 1668 644
rect 1602 -44 1668 68
rect 1760 644 1826 916
rect 1760 68 1766 644
rect 1820 68 1826 644
rect 1760 62 1826 68
rect 1918 644 1984 650
rect 1918 68 1924 644
rect 1978 68 1984 644
rect 1918 -44 1984 68
rect 2076 644 2142 916
rect 2076 68 2082 644
rect 2136 68 2142 644
rect 2076 62 2142 68
rect 2234 644 2300 650
rect 2234 68 2240 644
rect 2294 68 2300 644
rect 2234 -44 2300 68
rect 2392 644 2458 916
rect 2392 68 2398 644
rect 2452 68 2458 644
rect 2392 62 2458 68
rect 2860 60 3524 184
rect 256 -136 2300 -44
rect 2760 -38 2824 -32
rect 174 -414 240 -408
rect 174 -590 180 -414
rect 234 -590 240 -414
rect 174 -722 240 -590
rect 366 -414 432 -408
rect 366 -590 372 -414
rect 426 -590 432 -414
rect 366 -722 432 -590
rect 558 -414 624 -408
rect 558 -590 564 -414
rect 618 -590 624 -414
rect 558 -722 624 -590
rect 892 -414 956 -136
rect 892 -590 898 -414
rect 950 -590 956 -414
rect 892 -596 956 -590
rect 988 -414 1054 -408
rect 988 -590 994 -414
rect 1048 -590 1054 -414
rect 988 -722 1054 -590
rect 1086 -414 1150 -136
rect 1086 -590 1092 -414
rect 1144 -590 1150 -414
rect 1086 -596 1150 -590
rect 1182 -414 1248 -408
rect 1182 -590 1188 -414
rect 1240 -590 1248 -414
rect 1182 -722 1248 -590
rect 1278 -414 1342 -136
rect 1278 -590 1284 -414
rect 1336 -590 1342 -414
rect 1278 -596 1342 -590
rect 1374 -414 1438 -408
rect 1374 -590 1380 -414
rect 1432 -590 1438 -414
rect 1374 -722 1438 -590
rect 2760 -590 2766 -38
rect 2818 -590 2824 -38
rect 2760 -722 2824 -590
rect 2860 -38 2924 60
rect 2860 -590 2866 -38
rect 2918 -590 2924 -38
rect 2860 -596 2924 -590
rect 2956 -38 3020 -32
rect 2956 -590 2962 -38
rect 3014 -590 3020 -38
rect 2956 -722 3020 -590
rect 3052 -38 3116 60
rect 3052 -590 3058 -38
rect 3110 -590 3116 -38
rect 3052 -596 3116 -590
rect 3148 -38 3212 -32
rect 3148 -590 3154 -38
rect 3206 -590 3212 -38
rect 3148 -722 3212 -590
rect 3244 -38 3308 60
rect 3244 -590 3250 -38
rect 3302 -590 3308 -38
rect 3244 -596 3308 -590
rect 3400 -690 3524 60
rect 3584 -482 3590 936
rect 3642 -482 3648 936
rect 3714 936 3778 1068
rect 3714 -482 3720 936
rect 3772 -482 3778 936
rect 3844 936 3908 942
rect 3844 -482 3850 936
rect 3902 -482 3908 936
rect 3970 936 4034 1068
rect 3970 -482 3976 936
rect 4028 -482 4034 936
rect 4100 936 4164 942
rect 4100 -482 4106 936
rect 4158 -482 4164 936
rect 4226 936 4290 1068
rect 4226 -482 4232 936
rect 4284 -482 4290 936
rect 4356 936 4420 942
rect 4356 -482 4362 936
rect 4414 -482 4420 936
rect 4482 936 4546 1068
rect 4482 -482 4488 936
rect 4540 -482 4546 936
rect 4612 936 4676 942
rect 4612 -482 4618 936
rect 4670 -482 4676 936
rect 4738 936 4802 1068
rect 4738 -482 4744 936
rect 4796 -482 4802 936
rect 4868 936 4932 942
rect 4868 -482 4874 936
rect 4926 -482 4932 936
rect 4994 936 5058 1068
rect 4994 -482 5000 936
rect 5052 -482 5058 936
rect 5124 936 5188 942
rect 5124 -482 5130 936
rect 5182 -482 5188 936
rect 5250 936 5314 1068
rect 5250 -482 5256 936
rect 5308 -482 5314 936
rect 5380 936 5444 942
rect 5380 -482 5386 936
rect 5438 -482 5444 936
rect 5506 936 5570 1068
rect 5506 -482 5512 936
rect 5564 -482 5570 936
rect 3584 -690 3648 -482
rect 3844 -690 3908 -482
rect 4100 -690 4164 -482
rect 4356 -690 4420 -482
rect 4612 -690 4676 -482
rect 4868 -690 4932 -482
rect 5124 -690 5188 -482
rect 5380 -690 5444 -482
rect 174 -732 3290 -722
rect 174 -784 240 -732
rect 596 -784 994 -732
rect 1352 -734 3290 -732
rect 1352 -784 2818 -734
rect 174 -788 2818 -784
rect 3250 -788 3290 -734
rect 174 -812 3290 -788
rect 1618 -954 3272 -812
rect 3400 -814 5444 -690
rect 3560 -894 4734 -814
rect 3560 -1046 3570 -894
rect 4672 -1046 4734 -894
rect 3560 -1056 4734 -1046
<< via2 >>
rect 2922 1494 3386 1780
rect 3570 -1046 4672 -894
<< metal3 >>
rect 2912 1780 3396 1790
rect 2912 1570 2922 1780
rect 2878 1494 2922 1570
rect 3386 1570 3396 1780
rect 3386 1494 3428 1570
rect 2878 1222 3428 1494
rect 3560 -894 4680 -886
rect 3560 -1046 3570 -894
rect 4672 -1046 4680 -894
rect 3560 -1056 4680 -1046
<< via3 >>
rect 2922 1494 3386 1780
rect 3570 -1046 4672 -894
<< metal4 >>
rect 2910 1780 3396 1790
rect 2910 1494 2922 1780
rect 3386 1494 3396 1780
rect 2910 1484 3396 1494
rect 3560 -894 4680 -632
rect 3560 -1046 3570 -894
rect 4672 -1046 4680 -894
rect 3560 -1056 4680 -1046
<< via4 >>
rect 2922 1494 3386 1780
<< metal5 >>
rect 2878 1780 3428 1822
rect 2878 1494 2922 1780
rect 3386 1494 3428 1780
rect 2878 1222 3428 1494
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_0
timestamp 1665661446
transform -1 0 3767 0 -1 296
box -1150 -1100 1049 1100
use sky130_fd_pr__cap_mim_m3_2_6ZNTNB  sky130_fd_pr__cap_mim_m3_2_6ZNTNB_0
timestamp 1665661005
transform 1 0 4067 0 1 296
box -1351 -1100 849 1100
use sky130_fd_pr__nfet_01v8_lvt_46VND8  sky130_fd_pr__nfet_01v8_lvt_46VND8_0
timestamp 1665942972
transform 1 0 3035 0 1 -314
box -407 -498 407 498
use sky130_fd_pr__nfet_01v8_lvt_595QY5  sky130_fd_pr__nfet_01v8_lvt_595QY5_0
timestamp 1665942907
transform 1 0 351 0 1 -502
box -407 -310 407 310
use sky130_fd_pr__nfet_01v8_lvt_595QY5  sky130_fd_pr__nfet_01v8_lvt_595QY5_1
timestamp 1665942907
transform 1 0 1166 0 1 -502
box -407 -310 407 310
use sky130_fd_pr__nfet_03v3_nvt_QBNVYP  sky130_fd_pr__nfet_03v3_nvt_QBNVYP_0
timestamp 1665943141
transform 1 0 605 0 1 356
box -673 -558 673 558
use sky130_fd_pr__nfet_03v3_nvt_QBNVYP  sky130_fd_pr__nfet_03v3_nvt_QBNVYP_1
timestamp 1665943141
transform 1 0 1953 0 1 356
box -673 -558 673 558
use sky130_fd_pr__pfet_01v8_lvt_E98R26  sky130_fd_pr__pfet_01v8_lvt_E98R26_0
timestamp 1665943203
transform 1 0 183 0 1 1423
box -487 -507 487 507
use sky130_fd_pr__pfet_01v8_lvt_E98R26  sky130_fd_pr__pfet_01v8_lvt_E98R26_1
timestamp 1665943203
transform 1 0 1764 0 1 1423
box -487 -507 487 507
use sky130_fd_pr__pfet_01v8_lvt_ZUTRP2  sky130_fd_pr__pfet_01v8_lvt_ZUTRP2_0
timestamp 1665663699
transform 1 0 4579 0 1 227
box -1127 -939 1127 939
use sky130_fd_pr__res_xhigh_po_0p35_LSEQGR  sky130_fd_pr__res_xhigh_po_0p35_LSEQGR_0
timestamp 1665662444
transform 1 0 -259 0 1 -139
box -201 -673 201 673
<< labels >>
rlabel metal1 -446 -142 -446 -142 7 NonInv
port 2 w
rlabel metal2 2982 -930 2984 -930 5 Vss
port 5 s
rlabel metal2 2468 1216 2468 1216 1 Vdd
port 4 n
rlabel via3 3844 -950 3844 -950 5 Out
port 3 s
rlabel metal1 -456 -16 -456 -16 7 Inv
port 1 w
<< end >>
