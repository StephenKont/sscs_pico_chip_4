magic
tech sky130A
magscale 1 2
timestamp 1667067748
<< metal4 >>
rect -411 100750 -91 100800
rect -3351 97810 2849 100750
rect -3401 97490 2899 97810
rect -3351 94550 2849 97490
rect -411 94450 -91 94550
rect -3351 91510 2849 94450
rect -3401 91190 2899 91510
rect -3351 88250 2849 91190
rect -411 88150 -91 88250
rect -3351 85210 2849 88150
rect -3401 84890 2899 85210
rect -3351 81950 2849 84890
rect -411 81850 -91 81950
rect -3351 78910 2849 81850
rect -3401 78590 2899 78910
rect -3351 75650 2849 78590
rect -411 75550 -91 75650
rect -3351 72610 2849 75550
rect -3401 72290 2899 72610
rect -3351 69350 2849 72290
rect -411 69250 -91 69350
rect -3351 66310 2849 69250
rect -3401 65990 2899 66310
rect -3351 63050 2849 65990
rect -411 62950 -91 63050
rect -3351 60010 2849 62950
rect -3401 59690 2899 60010
rect -3351 56750 2849 59690
rect -411 56650 -91 56750
rect -3351 53710 2849 56650
rect -3401 53390 2899 53710
rect -3351 50450 2849 53390
rect -411 50350 -91 50450
rect -3351 47410 2849 50350
rect -3401 47090 2899 47410
rect -3351 44150 2849 47090
rect -411 44050 -91 44150
rect -3351 41110 2849 44050
rect -3401 40790 2899 41110
rect -3351 37850 2849 40790
rect -411 37750 -91 37850
rect -3351 34810 2849 37750
rect -3401 34490 2899 34810
rect -3351 31550 2849 34490
rect -411 31450 -91 31550
rect -3351 28510 2849 31450
rect -3401 28190 2899 28510
rect -3351 25250 2849 28190
rect -411 25150 -91 25250
rect -3351 22210 2849 25150
rect -3401 21890 2899 22210
rect -3351 18950 2849 21890
rect -411 18850 -91 18950
rect -3351 15910 2849 18850
rect -3401 15590 2899 15910
rect -3351 12650 2849 15590
rect -411 12550 -91 12650
rect -3351 9610 2849 12550
rect -3401 9290 2899 9610
rect -3351 6350 2849 9290
rect -411 6250 -91 6350
rect -3351 3310 2849 6250
rect -3401 2990 2899 3310
rect -3351 50 2849 2990
rect -411 -50 -91 50
rect -3351 -2990 2849 -50
rect -3401 -3310 2899 -2990
rect -3351 -6250 2849 -3310
rect -411 -6350 -91 -6250
rect -3351 -9290 2849 -6350
rect -3401 -9610 2899 -9290
rect -3351 -12550 2849 -9610
rect -411 -12650 -91 -12550
rect -3351 -15590 2849 -12650
rect -3401 -15910 2899 -15590
rect -3351 -18850 2849 -15910
rect -411 -18950 -91 -18850
rect -3351 -21890 2849 -18950
rect -3401 -22210 2899 -21890
rect -3351 -25150 2849 -22210
rect -411 -25250 -91 -25150
rect -3351 -28190 2849 -25250
rect -3401 -28510 2899 -28190
rect -3351 -31450 2849 -28510
rect -411 -31550 -91 -31450
rect -3351 -34490 2849 -31550
rect -3401 -34810 2899 -34490
rect -3351 -37750 2849 -34810
rect -411 -37850 -91 -37750
rect -3351 -40790 2849 -37850
rect -3401 -41110 2899 -40790
rect -3351 -44050 2849 -41110
rect -411 -44150 -91 -44050
rect -3351 -47090 2849 -44150
rect -3401 -47410 2899 -47090
rect -3351 -50350 2849 -47410
rect -411 -50450 -91 -50350
rect -3351 -53390 2849 -50450
rect -3401 -53710 2899 -53390
rect -3351 -56650 2849 -53710
rect -411 -56750 -91 -56650
rect -3351 -59690 2849 -56750
rect -3401 -60010 2899 -59690
rect -3351 -62950 2849 -60010
rect -411 -63050 -91 -62950
rect -3351 -65990 2849 -63050
rect -3401 -66310 2899 -65990
rect -3351 -69250 2849 -66310
rect -411 -69350 -91 -69250
rect -3351 -72290 2849 -69350
rect -3401 -72610 2899 -72290
rect -3351 -75550 2849 -72610
rect -411 -75650 -91 -75550
rect -3351 -78590 2849 -75650
rect -3401 -78910 2899 -78590
rect -3351 -81850 2849 -78910
rect -411 -81950 -91 -81850
rect -3351 -84890 2849 -81950
rect -3401 -85210 2899 -84890
rect -3351 -88150 2849 -85210
rect -411 -88250 -91 -88150
rect -3351 -91190 2849 -88250
rect -3401 -91510 2899 -91190
rect -3351 -94450 2849 -91510
rect -411 -94550 -91 -94450
rect -3351 -97490 2849 -94550
rect -3401 -97810 2899 -97490
rect -3351 -100750 2849 -97810
rect -411 -100800 -91 -100750
<< mimcap2 >>
rect -3251 100610 2749 100650
rect -3251 94690 -3211 100610
rect 2625 94690 2749 100610
rect -3251 94650 2749 94690
rect -3251 94310 2749 94350
rect -3251 88390 -3211 94310
rect 2625 88390 2749 94310
rect -3251 88350 2749 88390
rect -3251 88010 2749 88050
rect -3251 82090 -3211 88010
rect 2625 82090 2749 88010
rect -3251 82050 2749 82090
rect -3251 81710 2749 81750
rect -3251 75790 -3211 81710
rect 2625 75790 2749 81710
rect -3251 75750 2749 75790
rect -3251 75410 2749 75450
rect -3251 69490 -3211 75410
rect 2625 69490 2749 75410
rect -3251 69450 2749 69490
rect -3251 69110 2749 69150
rect -3251 63190 -3211 69110
rect 2625 63190 2749 69110
rect -3251 63150 2749 63190
rect -3251 62810 2749 62850
rect -3251 56890 -3211 62810
rect 2625 56890 2749 62810
rect -3251 56850 2749 56890
rect -3251 56510 2749 56550
rect -3251 50590 -3211 56510
rect 2625 50590 2749 56510
rect -3251 50550 2749 50590
rect -3251 50210 2749 50250
rect -3251 44290 -3211 50210
rect 2625 44290 2749 50210
rect -3251 44250 2749 44290
rect -3251 43910 2749 43950
rect -3251 37990 -3211 43910
rect 2625 37990 2749 43910
rect -3251 37950 2749 37990
rect -3251 37610 2749 37650
rect -3251 31690 -3211 37610
rect 2625 31690 2749 37610
rect -3251 31650 2749 31690
rect -3251 31310 2749 31350
rect -3251 25390 -3211 31310
rect 2625 25390 2749 31310
rect -3251 25350 2749 25390
rect -3251 25010 2749 25050
rect -3251 19090 -3211 25010
rect 2625 19090 2749 25010
rect -3251 19050 2749 19090
rect -3251 18710 2749 18750
rect -3251 12790 -3211 18710
rect 2625 12790 2749 18710
rect -3251 12750 2749 12790
rect -3251 12410 2749 12450
rect -3251 6490 -3211 12410
rect 2625 6490 2749 12410
rect -3251 6450 2749 6490
rect -3251 6110 2749 6150
rect -3251 190 -3211 6110
rect 2625 190 2749 6110
rect -3251 150 2749 190
rect -3251 -190 2749 -150
rect -3251 -6110 -3211 -190
rect 2625 -6110 2749 -190
rect -3251 -6150 2749 -6110
rect -3251 -6490 2749 -6450
rect -3251 -12410 -3211 -6490
rect 2625 -12410 2749 -6490
rect -3251 -12450 2749 -12410
rect -3251 -12790 2749 -12750
rect -3251 -18710 -3211 -12790
rect 2625 -18710 2749 -12790
rect -3251 -18750 2749 -18710
rect -3251 -19090 2749 -19050
rect -3251 -25010 -3211 -19090
rect 2625 -25010 2749 -19090
rect -3251 -25050 2749 -25010
rect -3251 -25390 2749 -25350
rect -3251 -31310 -3211 -25390
rect 2625 -31310 2749 -25390
rect -3251 -31350 2749 -31310
rect -3251 -31690 2749 -31650
rect -3251 -37610 -3211 -31690
rect 2625 -37610 2749 -31690
rect -3251 -37650 2749 -37610
rect -3251 -37990 2749 -37950
rect -3251 -43910 -3211 -37990
rect 2625 -43910 2749 -37990
rect -3251 -43950 2749 -43910
rect -3251 -44290 2749 -44250
rect -3251 -50210 -3211 -44290
rect 2625 -50210 2749 -44290
rect -3251 -50250 2749 -50210
rect -3251 -50590 2749 -50550
rect -3251 -56510 -3211 -50590
rect 2625 -56510 2749 -50590
rect -3251 -56550 2749 -56510
rect -3251 -56890 2749 -56850
rect -3251 -62810 -3211 -56890
rect 2625 -62810 2749 -56890
rect -3251 -62850 2749 -62810
rect -3251 -63190 2749 -63150
rect -3251 -69110 -3211 -63190
rect 2625 -69110 2749 -63190
rect -3251 -69150 2749 -69110
rect -3251 -69490 2749 -69450
rect -3251 -75410 -3211 -69490
rect 2625 -75410 2749 -69490
rect -3251 -75450 2749 -75410
rect -3251 -75790 2749 -75750
rect -3251 -81710 -3211 -75790
rect 2625 -81710 2749 -75790
rect -3251 -81750 2749 -81710
rect -3251 -82090 2749 -82050
rect -3251 -88010 -3211 -82090
rect 2625 -88010 2749 -82090
rect -3251 -88050 2749 -88010
rect -3251 -88390 2749 -88350
rect -3251 -94310 -3211 -88390
rect 2625 -94310 2749 -88390
rect -3251 -94350 2749 -94310
rect -3251 -94690 2749 -94650
rect -3251 -100610 -3211 -94690
rect 2625 -100610 2749 -94690
rect -3251 -100650 2749 -100610
<< mimcap2contact >>
rect -3211 94690 2625 100610
rect -3211 88390 2625 94310
rect -3211 82090 2625 88010
rect -3211 75790 2625 81710
rect -3211 69490 2625 75410
rect -3211 63190 2625 69110
rect -3211 56890 2625 62810
rect -3211 50590 2625 56510
rect -3211 44290 2625 50210
rect -3211 37990 2625 43910
rect -3211 31690 2625 37610
rect -3211 25390 2625 31310
rect -3211 19090 2625 25010
rect -3211 12790 2625 18710
rect -3211 6490 2625 12410
rect -3211 190 2625 6110
rect -3211 -6110 2625 -190
rect -3211 -12410 2625 -6490
rect -3211 -18710 2625 -12790
rect -3211 -25010 2625 -19090
rect -3211 -31310 2625 -25390
rect -3211 -37610 2625 -31690
rect -3211 -43910 2625 -37990
rect -3211 -50210 2625 -44290
rect -3211 -56510 2625 -50590
rect -3211 -62810 2625 -56890
rect -3211 -69110 2625 -63190
rect -3211 -75410 2625 -69490
rect -3211 -81710 2625 -75790
rect -3211 -88010 2625 -82090
rect -3211 -94310 2625 -88390
rect -3211 -100610 2625 -94690
<< metal5 >>
rect -411 100634 -91 100800
rect -3235 100610 2649 100634
rect -3235 97810 -3211 100610
rect -3401 97490 -3211 97810
rect -3235 94690 -3211 97490
rect 2625 97810 2649 100610
rect 2625 97490 2899 97810
rect 2625 94690 2649 97490
rect -3235 94666 2649 94690
rect -411 94334 -91 94666
rect -3235 94310 2649 94334
rect -3235 91510 -3211 94310
rect -3401 91190 -3211 91510
rect -3235 88390 -3211 91190
rect 2625 91510 2649 94310
rect 2625 91190 2899 91510
rect 2625 88390 2649 91190
rect -3235 88366 2649 88390
rect -411 88034 -91 88366
rect -3235 88010 2649 88034
rect -3235 85210 -3211 88010
rect -3401 84890 -3211 85210
rect -3235 82090 -3211 84890
rect 2625 85210 2649 88010
rect 2625 84890 2899 85210
rect 2625 82090 2649 84890
rect -3235 82066 2649 82090
rect -411 81734 -91 82066
rect -3235 81710 2649 81734
rect -3235 78910 -3211 81710
rect -3401 78590 -3211 78910
rect -3235 75790 -3211 78590
rect 2625 78910 2649 81710
rect 2625 78590 2899 78910
rect 2625 75790 2649 78590
rect -3235 75766 2649 75790
rect -411 75434 -91 75766
rect -3235 75410 2649 75434
rect -3235 72610 -3211 75410
rect -3401 72290 -3211 72610
rect -3235 69490 -3211 72290
rect 2625 72610 2649 75410
rect 2625 72290 2899 72610
rect 2625 69490 2649 72290
rect -3235 69466 2649 69490
rect -411 69134 -91 69466
rect -3235 69110 2649 69134
rect -3235 66310 -3211 69110
rect -3401 65990 -3211 66310
rect -3235 63190 -3211 65990
rect 2625 66310 2649 69110
rect 2625 65990 2899 66310
rect 2625 63190 2649 65990
rect -3235 63166 2649 63190
rect -411 62834 -91 63166
rect -3235 62810 2649 62834
rect -3235 60010 -3211 62810
rect -3401 59690 -3211 60010
rect -3235 56890 -3211 59690
rect 2625 60010 2649 62810
rect 2625 59690 2899 60010
rect 2625 56890 2649 59690
rect -3235 56866 2649 56890
rect -411 56534 -91 56866
rect -3235 56510 2649 56534
rect -3235 53710 -3211 56510
rect -3401 53390 -3211 53710
rect -3235 50590 -3211 53390
rect 2625 53710 2649 56510
rect 2625 53390 2899 53710
rect 2625 50590 2649 53390
rect -3235 50566 2649 50590
rect -411 50234 -91 50566
rect -3235 50210 2649 50234
rect -3235 47410 -3211 50210
rect -3401 47090 -3211 47410
rect -3235 44290 -3211 47090
rect 2625 47410 2649 50210
rect 2625 47090 2899 47410
rect 2625 44290 2649 47090
rect -3235 44266 2649 44290
rect -411 43934 -91 44266
rect -3235 43910 2649 43934
rect -3235 41110 -3211 43910
rect -3401 40790 -3211 41110
rect -3235 37990 -3211 40790
rect 2625 41110 2649 43910
rect 2625 40790 2899 41110
rect 2625 37990 2649 40790
rect -3235 37966 2649 37990
rect -411 37634 -91 37966
rect -3235 37610 2649 37634
rect -3235 34810 -3211 37610
rect -3401 34490 -3211 34810
rect -3235 31690 -3211 34490
rect 2625 34810 2649 37610
rect 2625 34490 2899 34810
rect 2625 31690 2649 34490
rect -3235 31666 2649 31690
rect -411 31334 -91 31666
rect -3235 31310 2649 31334
rect -3235 28510 -3211 31310
rect -3401 28190 -3211 28510
rect -3235 25390 -3211 28190
rect 2625 28510 2649 31310
rect 2625 28190 2899 28510
rect 2625 25390 2649 28190
rect -3235 25366 2649 25390
rect -411 25034 -91 25366
rect -3235 25010 2649 25034
rect -3235 22210 -3211 25010
rect -3401 21890 -3211 22210
rect -3235 19090 -3211 21890
rect 2625 22210 2649 25010
rect 2625 21890 2899 22210
rect 2625 19090 2649 21890
rect -3235 19066 2649 19090
rect -411 18734 -91 19066
rect -3235 18710 2649 18734
rect -3235 15910 -3211 18710
rect -3401 15590 -3211 15910
rect -3235 12790 -3211 15590
rect 2625 15910 2649 18710
rect 2625 15590 2899 15910
rect 2625 12790 2649 15590
rect -3235 12766 2649 12790
rect -411 12434 -91 12766
rect -3235 12410 2649 12434
rect -3235 9610 -3211 12410
rect -3401 9290 -3211 9610
rect -3235 6490 -3211 9290
rect 2625 9610 2649 12410
rect 2625 9290 2899 9610
rect 2625 6490 2649 9290
rect -3235 6466 2649 6490
rect -411 6134 -91 6466
rect -3235 6110 2649 6134
rect -3235 3310 -3211 6110
rect -3401 2990 -3211 3310
rect -3235 190 -3211 2990
rect 2625 3310 2649 6110
rect 2625 2990 2899 3310
rect 2625 190 2649 2990
rect -3235 166 2649 190
rect -411 -166 -91 166
rect -3235 -190 2649 -166
rect -3235 -2990 -3211 -190
rect -3401 -3310 -3211 -2990
rect -3235 -6110 -3211 -3310
rect 2625 -2990 2649 -190
rect 2625 -3310 2899 -2990
rect 2625 -6110 2649 -3310
rect -3235 -6134 2649 -6110
rect -411 -6466 -91 -6134
rect -3235 -6490 2649 -6466
rect -3235 -9290 -3211 -6490
rect -3401 -9610 -3211 -9290
rect -3235 -12410 -3211 -9610
rect 2625 -9290 2649 -6490
rect 2625 -9610 2899 -9290
rect 2625 -12410 2649 -9610
rect -3235 -12434 2649 -12410
rect -411 -12766 -91 -12434
rect -3235 -12790 2649 -12766
rect -3235 -15590 -3211 -12790
rect -3401 -15910 -3211 -15590
rect -3235 -18710 -3211 -15910
rect 2625 -15590 2649 -12790
rect 2625 -15910 2899 -15590
rect 2625 -18710 2649 -15910
rect -3235 -18734 2649 -18710
rect -411 -19066 -91 -18734
rect -3235 -19090 2649 -19066
rect -3235 -21890 -3211 -19090
rect -3401 -22210 -3211 -21890
rect -3235 -25010 -3211 -22210
rect 2625 -21890 2649 -19090
rect 2625 -22210 2899 -21890
rect 2625 -25010 2649 -22210
rect -3235 -25034 2649 -25010
rect -411 -25366 -91 -25034
rect -3235 -25390 2649 -25366
rect -3235 -28190 -3211 -25390
rect -3401 -28510 -3211 -28190
rect -3235 -31310 -3211 -28510
rect 2625 -28190 2649 -25390
rect 2625 -28510 2899 -28190
rect 2625 -31310 2649 -28510
rect -3235 -31334 2649 -31310
rect -411 -31666 -91 -31334
rect -3235 -31690 2649 -31666
rect -3235 -34490 -3211 -31690
rect -3401 -34810 -3211 -34490
rect -3235 -37610 -3211 -34810
rect 2625 -34490 2649 -31690
rect 2625 -34810 2899 -34490
rect 2625 -37610 2649 -34810
rect -3235 -37634 2649 -37610
rect -411 -37966 -91 -37634
rect -3235 -37990 2649 -37966
rect -3235 -40790 -3211 -37990
rect -3401 -41110 -3211 -40790
rect -3235 -43910 -3211 -41110
rect 2625 -40790 2649 -37990
rect 2625 -41110 2899 -40790
rect 2625 -43910 2649 -41110
rect -3235 -43934 2649 -43910
rect -411 -44266 -91 -43934
rect -3235 -44290 2649 -44266
rect -3235 -47090 -3211 -44290
rect -3401 -47410 -3211 -47090
rect -3235 -50210 -3211 -47410
rect 2625 -47090 2649 -44290
rect 2625 -47410 2899 -47090
rect 2625 -50210 2649 -47410
rect -3235 -50234 2649 -50210
rect -411 -50566 -91 -50234
rect -3235 -50590 2649 -50566
rect -3235 -53390 -3211 -50590
rect -3401 -53710 -3211 -53390
rect -3235 -56510 -3211 -53710
rect 2625 -53390 2649 -50590
rect 2625 -53710 2899 -53390
rect 2625 -56510 2649 -53710
rect -3235 -56534 2649 -56510
rect -411 -56866 -91 -56534
rect -3235 -56890 2649 -56866
rect -3235 -59690 -3211 -56890
rect -3401 -60010 -3211 -59690
rect -3235 -62810 -3211 -60010
rect 2625 -59690 2649 -56890
rect 2625 -60010 2899 -59690
rect 2625 -62810 2649 -60010
rect -3235 -62834 2649 -62810
rect -411 -63166 -91 -62834
rect -3235 -63190 2649 -63166
rect -3235 -65990 -3211 -63190
rect -3401 -66310 -3211 -65990
rect -3235 -69110 -3211 -66310
rect 2625 -65990 2649 -63190
rect 2625 -66310 2899 -65990
rect 2625 -69110 2649 -66310
rect -3235 -69134 2649 -69110
rect -411 -69466 -91 -69134
rect -3235 -69490 2649 -69466
rect -3235 -72290 -3211 -69490
rect -3401 -72610 -3211 -72290
rect -3235 -75410 -3211 -72610
rect 2625 -72290 2649 -69490
rect 2625 -72610 2899 -72290
rect 2625 -75410 2649 -72610
rect -3235 -75434 2649 -75410
rect -411 -75766 -91 -75434
rect -3235 -75790 2649 -75766
rect -3235 -78590 -3211 -75790
rect -3401 -78910 -3211 -78590
rect -3235 -81710 -3211 -78910
rect 2625 -78590 2649 -75790
rect 2625 -78910 2899 -78590
rect 2625 -81710 2649 -78910
rect -3235 -81734 2649 -81710
rect -411 -82066 -91 -81734
rect -3235 -82090 2649 -82066
rect -3235 -84890 -3211 -82090
rect -3401 -85210 -3211 -84890
rect -3235 -88010 -3211 -85210
rect 2625 -84890 2649 -82090
rect 2625 -85210 2899 -84890
rect 2625 -88010 2649 -85210
rect -3235 -88034 2649 -88010
rect -411 -88366 -91 -88034
rect -3235 -88390 2649 -88366
rect -3235 -91190 -3211 -88390
rect -3401 -91510 -3211 -91190
rect -3235 -94310 -3211 -91510
rect 2625 -91190 2649 -88390
rect 2625 -91510 2899 -91190
rect 2625 -94310 2649 -91510
rect -3235 -94334 2649 -94310
rect -411 -94666 -91 -94334
rect -3235 -94690 2649 -94666
rect -3235 -97490 -3211 -94690
rect -3401 -97810 -3211 -97490
rect -3235 -100610 -3211 -97810
rect 2625 -97490 2649 -94690
rect 2625 -97810 2899 -97490
rect 2625 -100610 2649 -97810
rect -3235 -100634 2649 -100610
rect -411 -100800 -91 -100634
<< properties >>
string FIXED_BBOX -3351 94550 2849 100750
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 32 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
