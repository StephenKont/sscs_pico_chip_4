magic
tech sky130A
magscale 1 2
timestamp 1665560597
<< nwell >>
rect -358 -4193 358 4193
<< mvpmos >>
rect -100 3496 100 3896
rect -100 2968 100 3368
rect -100 2440 100 2840
rect -100 1912 100 2312
rect -100 1384 100 1784
rect -100 856 100 1256
rect -100 328 100 728
rect -100 -200 100 200
rect -100 -728 100 -328
rect -100 -1256 100 -856
rect -100 -1784 100 -1384
rect -100 -2312 100 -1912
rect -100 -2840 100 -2440
rect -100 -3368 100 -2968
rect -100 -3896 100 -3496
<< mvpdiff >>
rect -158 3884 -100 3896
rect -158 3508 -146 3884
rect -112 3508 -100 3884
rect -158 3496 -100 3508
rect 100 3884 158 3896
rect 100 3508 112 3884
rect 146 3508 158 3884
rect 100 3496 158 3508
rect -158 3356 -100 3368
rect -158 2980 -146 3356
rect -112 2980 -100 3356
rect -158 2968 -100 2980
rect 100 3356 158 3368
rect 100 2980 112 3356
rect 146 2980 158 3356
rect 100 2968 158 2980
rect -158 2828 -100 2840
rect -158 2452 -146 2828
rect -112 2452 -100 2828
rect -158 2440 -100 2452
rect 100 2828 158 2840
rect 100 2452 112 2828
rect 146 2452 158 2828
rect 100 2440 158 2452
rect -158 2300 -100 2312
rect -158 1924 -146 2300
rect -112 1924 -100 2300
rect -158 1912 -100 1924
rect 100 2300 158 2312
rect 100 1924 112 2300
rect 146 1924 158 2300
rect 100 1912 158 1924
rect -158 1772 -100 1784
rect -158 1396 -146 1772
rect -112 1396 -100 1772
rect -158 1384 -100 1396
rect 100 1772 158 1784
rect 100 1396 112 1772
rect 146 1396 158 1772
rect 100 1384 158 1396
rect -158 1244 -100 1256
rect -158 868 -146 1244
rect -112 868 -100 1244
rect -158 856 -100 868
rect 100 1244 158 1256
rect 100 868 112 1244
rect 146 868 158 1244
rect 100 856 158 868
rect -158 716 -100 728
rect -158 340 -146 716
rect -112 340 -100 716
rect -158 328 -100 340
rect 100 716 158 728
rect 100 340 112 716
rect 146 340 158 716
rect 100 328 158 340
rect -158 188 -100 200
rect -158 -188 -146 188
rect -112 -188 -100 188
rect -158 -200 -100 -188
rect 100 188 158 200
rect 100 -188 112 188
rect 146 -188 158 188
rect 100 -200 158 -188
rect -158 -340 -100 -328
rect -158 -716 -146 -340
rect -112 -716 -100 -340
rect -158 -728 -100 -716
rect 100 -340 158 -328
rect 100 -716 112 -340
rect 146 -716 158 -340
rect 100 -728 158 -716
rect -158 -868 -100 -856
rect -158 -1244 -146 -868
rect -112 -1244 -100 -868
rect -158 -1256 -100 -1244
rect 100 -868 158 -856
rect 100 -1244 112 -868
rect 146 -1244 158 -868
rect 100 -1256 158 -1244
rect -158 -1396 -100 -1384
rect -158 -1772 -146 -1396
rect -112 -1772 -100 -1396
rect -158 -1784 -100 -1772
rect 100 -1396 158 -1384
rect 100 -1772 112 -1396
rect 146 -1772 158 -1396
rect 100 -1784 158 -1772
rect -158 -1924 -100 -1912
rect -158 -2300 -146 -1924
rect -112 -2300 -100 -1924
rect -158 -2312 -100 -2300
rect 100 -1924 158 -1912
rect 100 -2300 112 -1924
rect 146 -2300 158 -1924
rect 100 -2312 158 -2300
rect -158 -2452 -100 -2440
rect -158 -2828 -146 -2452
rect -112 -2828 -100 -2452
rect -158 -2840 -100 -2828
rect 100 -2452 158 -2440
rect 100 -2828 112 -2452
rect 146 -2828 158 -2452
rect 100 -2840 158 -2828
rect -158 -2980 -100 -2968
rect -158 -3356 -146 -2980
rect -112 -3356 -100 -2980
rect -158 -3368 -100 -3356
rect 100 -2980 158 -2968
rect 100 -3356 112 -2980
rect 146 -3356 158 -2980
rect 100 -3368 158 -3356
rect -158 -3508 -100 -3496
rect -158 -3884 -146 -3508
rect -112 -3884 -100 -3508
rect -158 -3896 -100 -3884
rect 100 -3508 158 -3496
rect 100 -3884 112 -3508
rect 146 -3884 158 -3508
rect 100 -3896 158 -3884
<< mvpdiffc >>
rect -146 3508 -112 3884
rect 112 3508 146 3884
rect -146 2980 -112 3356
rect 112 2980 146 3356
rect -146 2452 -112 2828
rect 112 2452 146 2828
rect -146 1924 -112 2300
rect 112 1924 146 2300
rect -146 1396 -112 1772
rect 112 1396 146 1772
rect -146 868 -112 1244
rect 112 868 146 1244
rect -146 340 -112 716
rect 112 340 146 716
rect -146 -188 -112 188
rect 112 -188 146 188
rect -146 -716 -112 -340
rect 112 -716 146 -340
rect -146 -1244 -112 -868
rect 112 -1244 146 -868
rect -146 -1772 -112 -1396
rect 112 -1772 146 -1396
rect -146 -2300 -112 -1924
rect 112 -2300 146 -1924
rect -146 -2828 -112 -2452
rect 112 -2828 146 -2452
rect -146 -3356 -112 -2980
rect 112 -3356 146 -2980
rect -146 -3884 -112 -3508
rect 112 -3884 146 -3508
<< mvnsubdiff >>
rect -292 4115 292 4127
rect -292 4081 -184 4115
rect 184 4081 292 4115
rect -292 4069 292 4081
rect -292 4019 -234 4069
rect -292 -4019 -280 4019
rect -246 -4019 -234 4019
rect 234 4019 292 4069
rect -292 -4069 -234 -4019
rect 234 -4019 246 4019
rect 280 -4019 292 4019
rect 234 -4069 292 -4019
rect -292 -4081 292 -4069
rect -292 -4115 -184 -4081
rect 184 -4115 292 -4081
rect -292 -4127 292 -4115
<< mvnsubdiffcont >>
rect -184 4081 184 4115
rect -280 -4019 -246 4019
rect 246 -4019 280 4019
rect -184 -4115 184 -4081
<< poly >>
rect -100 3977 100 3993
rect -100 3943 -84 3977
rect 84 3943 100 3977
rect -100 3896 100 3943
rect -100 3449 100 3496
rect -100 3415 -84 3449
rect 84 3415 100 3449
rect -100 3368 100 3415
rect -100 2921 100 2968
rect -100 2887 -84 2921
rect 84 2887 100 2921
rect -100 2840 100 2887
rect -100 2393 100 2440
rect -100 2359 -84 2393
rect 84 2359 100 2393
rect -100 2312 100 2359
rect -100 1865 100 1912
rect -100 1831 -84 1865
rect 84 1831 100 1865
rect -100 1784 100 1831
rect -100 1337 100 1384
rect -100 1303 -84 1337
rect 84 1303 100 1337
rect -100 1256 100 1303
rect -100 809 100 856
rect -100 775 -84 809
rect 84 775 100 809
rect -100 728 100 775
rect -100 281 100 328
rect -100 247 -84 281
rect 84 247 100 281
rect -100 200 100 247
rect -100 -247 100 -200
rect -100 -281 -84 -247
rect 84 -281 100 -247
rect -100 -328 100 -281
rect -100 -775 100 -728
rect -100 -809 -84 -775
rect 84 -809 100 -775
rect -100 -856 100 -809
rect -100 -1303 100 -1256
rect -100 -1337 -84 -1303
rect 84 -1337 100 -1303
rect -100 -1384 100 -1337
rect -100 -1831 100 -1784
rect -100 -1865 -84 -1831
rect 84 -1865 100 -1831
rect -100 -1912 100 -1865
rect -100 -2359 100 -2312
rect -100 -2393 -84 -2359
rect 84 -2393 100 -2359
rect -100 -2440 100 -2393
rect -100 -2887 100 -2840
rect -100 -2921 -84 -2887
rect 84 -2921 100 -2887
rect -100 -2968 100 -2921
rect -100 -3415 100 -3368
rect -100 -3449 -84 -3415
rect 84 -3449 100 -3415
rect -100 -3496 100 -3449
rect -100 -3943 100 -3896
rect -100 -3977 -84 -3943
rect 84 -3977 100 -3943
rect -100 -3993 100 -3977
<< polycont >>
rect -84 3943 84 3977
rect -84 3415 84 3449
rect -84 2887 84 2921
rect -84 2359 84 2393
rect -84 1831 84 1865
rect -84 1303 84 1337
rect -84 775 84 809
rect -84 247 84 281
rect -84 -281 84 -247
rect -84 -809 84 -775
rect -84 -1337 84 -1303
rect -84 -1865 84 -1831
rect -84 -2393 84 -2359
rect -84 -2921 84 -2887
rect -84 -3449 84 -3415
rect -84 -3977 84 -3943
<< locali >>
rect -280 4081 -184 4115
rect 184 4081 280 4115
rect -280 4019 -246 4081
rect 246 4019 280 4081
rect -100 3943 -84 3977
rect 84 3943 100 3977
rect -146 3884 -112 3900
rect -146 3492 -112 3508
rect 112 3884 146 3900
rect 112 3492 146 3508
rect -100 3415 -84 3449
rect 84 3415 100 3449
rect -146 3356 -112 3372
rect -146 2964 -112 2980
rect 112 3356 146 3372
rect 112 2964 146 2980
rect -100 2887 -84 2921
rect 84 2887 100 2921
rect -146 2828 -112 2844
rect -146 2436 -112 2452
rect 112 2828 146 2844
rect 112 2436 146 2452
rect -100 2359 -84 2393
rect 84 2359 100 2393
rect -146 2300 -112 2316
rect -146 1908 -112 1924
rect 112 2300 146 2316
rect 112 1908 146 1924
rect -100 1831 -84 1865
rect 84 1831 100 1865
rect -146 1772 -112 1788
rect -146 1380 -112 1396
rect 112 1772 146 1788
rect 112 1380 146 1396
rect -100 1303 -84 1337
rect 84 1303 100 1337
rect -146 1244 -112 1260
rect -146 852 -112 868
rect 112 1244 146 1260
rect 112 852 146 868
rect -100 775 -84 809
rect 84 775 100 809
rect -146 716 -112 732
rect -146 324 -112 340
rect 112 716 146 732
rect 112 324 146 340
rect -100 247 -84 281
rect 84 247 100 281
rect -146 188 -112 204
rect -146 -204 -112 -188
rect 112 188 146 204
rect 112 -204 146 -188
rect -100 -281 -84 -247
rect 84 -281 100 -247
rect -146 -340 -112 -324
rect -146 -732 -112 -716
rect 112 -340 146 -324
rect 112 -732 146 -716
rect -100 -809 -84 -775
rect 84 -809 100 -775
rect -146 -868 -112 -852
rect -146 -1260 -112 -1244
rect 112 -868 146 -852
rect 112 -1260 146 -1244
rect -100 -1337 -84 -1303
rect 84 -1337 100 -1303
rect -146 -1396 -112 -1380
rect -146 -1788 -112 -1772
rect 112 -1396 146 -1380
rect 112 -1788 146 -1772
rect -100 -1865 -84 -1831
rect 84 -1865 100 -1831
rect -146 -1924 -112 -1908
rect -146 -2316 -112 -2300
rect 112 -1924 146 -1908
rect 112 -2316 146 -2300
rect -100 -2393 -84 -2359
rect 84 -2393 100 -2359
rect -146 -2452 -112 -2436
rect -146 -2844 -112 -2828
rect 112 -2452 146 -2436
rect 112 -2844 146 -2828
rect -100 -2921 -84 -2887
rect 84 -2921 100 -2887
rect -146 -2980 -112 -2964
rect -146 -3372 -112 -3356
rect 112 -2980 146 -2964
rect 112 -3372 146 -3356
rect -100 -3449 -84 -3415
rect 84 -3449 100 -3415
rect -146 -3508 -112 -3492
rect -146 -3900 -112 -3884
rect 112 -3508 146 -3492
rect 112 -3900 146 -3884
rect -100 -3977 -84 -3943
rect 84 -3977 100 -3943
rect -280 -4081 -246 -4019
rect 246 -4081 280 -4019
rect -280 -4115 -184 -4081
rect 184 -4115 280 -4081
<< viali >>
rect -84 3943 84 3977
rect -146 3508 -112 3884
rect 112 3508 146 3884
rect -84 3415 84 3449
rect -146 2980 -112 3356
rect 112 2980 146 3356
rect -84 2887 84 2921
rect -146 2452 -112 2828
rect 112 2452 146 2828
rect -84 2359 84 2393
rect -146 1924 -112 2300
rect 112 1924 146 2300
rect -84 1831 84 1865
rect -146 1396 -112 1772
rect 112 1396 146 1772
rect -84 1303 84 1337
rect -146 868 -112 1244
rect 112 868 146 1244
rect -84 775 84 809
rect -146 340 -112 716
rect 112 340 146 716
rect -84 247 84 281
rect -146 -188 -112 188
rect 112 -188 146 188
rect -84 -281 84 -247
rect -146 -716 -112 -340
rect 112 -716 146 -340
rect -84 -809 84 -775
rect -146 -1244 -112 -868
rect 112 -1244 146 -868
rect -84 -1337 84 -1303
rect -146 -1772 -112 -1396
rect 112 -1772 146 -1396
rect -84 -1865 84 -1831
rect -146 -2300 -112 -1924
rect 112 -2300 146 -1924
rect -84 -2393 84 -2359
rect -146 -2828 -112 -2452
rect 112 -2828 146 -2452
rect -84 -2921 84 -2887
rect -146 -3356 -112 -2980
rect 112 -3356 146 -2980
rect -84 -3449 84 -3415
rect -146 -3884 -112 -3508
rect 112 -3884 146 -3508
rect -84 -3977 84 -3943
<< metal1 >>
rect -96 3977 96 3983
rect -96 3943 -84 3977
rect 84 3943 96 3977
rect -96 3937 96 3943
rect -152 3884 -106 3896
rect -152 3508 -146 3884
rect -112 3508 -106 3884
rect -152 3496 -106 3508
rect 106 3884 152 3896
rect 106 3508 112 3884
rect 146 3508 152 3884
rect 106 3496 152 3508
rect -96 3449 96 3455
rect -96 3415 -84 3449
rect 84 3415 96 3449
rect -96 3409 96 3415
rect -152 3356 -106 3368
rect -152 2980 -146 3356
rect -112 2980 -106 3356
rect -152 2968 -106 2980
rect 106 3356 152 3368
rect 106 2980 112 3356
rect 146 2980 152 3356
rect 106 2968 152 2980
rect -96 2921 96 2927
rect -96 2887 -84 2921
rect 84 2887 96 2921
rect -96 2881 96 2887
rect -152 2828 -106 2840
rect -152 2452 -146 2828
rect -112 2452 -106 2828
rect -152 2440 -106 2452
rect 106 2828 152 2840
rect 106 2452 112 2828
rect 146 2452 152 2828
rect 106 2440 152 2452
rect -96 2393 96 2399
rect -96 2359 -84 2393
rect 84 2359 96 2393
rect -96 2353 96 2359
rect -152 2300 -106 2312
rect -152 1924 -146 2300
rect -112 1924 -106 2300
rect -152 1912 -106 1924
rect 106 2300 152 2312
rect 106 1924 112 2300
rect 146 1924 152 2300
rect 106 1912 152 1924
rect -96 1865 96 1871
rect -96 1831 -84 1865
rect 84 1831 96 1865
rect -96 1825 96 1831
rect -152 1772 -106 1784
rect -152 1396 -146 1772
rect -112 1396 -106 1772
rect -152 1384 -106 1396
rect 106 1772 152 1784
rect 106 1396 112 1772
rect 146 1396 152 1772
rect 106 1384 152 1396
rect -96 1337 96 1343
rect -96 1303 -84 1337
rect 84 1303 96 1337
rect -96 1297 96 1303
rect -152 1244 -106 1256
rect -152 868 -146 1244
rect -112 868 -106 1244
rect -152 856 -106 868
rect 106 1244 152 1256
rect 106 868 112 1244
rect 146 868 152 1244
rect 106 856 152 868
rect -96 809 96 815
rect -96 775 -84 809
rect 84 775 96 809
rect -96 769 96 775
rect -152 716 -106 728
rect -152 340 -146 716
rect -112 340 -106 716
rect -152 328 -106 340
rect 106 716 152 728
rect 106 340 112 716
rect 146 340 152 716
rect 106 328 152 340
rect -96 281 96 287
rect -96 247 -84 281
rect 84 247 96 281
rect -96 241 96 247
rect -152 188 -106 200
rect -152 -188 -146 188
rect -112 -188 -106 188
rect -152 -200 -106 -188
rect 106 188 152 200
rect 106 -188 112 188
rect 146 -188 152 188
rect 106 -200 152 -188
rect -96 -247 96 -241
rect -96 -281 -84 -247
rect 84 -281 96 -247
rect -96 -287 96 -281
rect -152 -340 -106 -328
rect -152 -716 -146 -340
rect -112 -716 -106 -340
rect -152 -728 -106 -716
rect 106 -340 152 -328
rect 106 -716 112 -340
rect 146 -716 152 -340
rect 106 -728 152 -716
rect -96 -775 96 -769
rect -96 -809 -84 -775
rect 84 -809 96 -775
rect -96 -815 96 -809
rect -152 -868 -106 -856
rect -152 -1244 -146 -868
rect -112 -1244 -106 -868
rect -152 -1256 -106 -1244
rect 106 -868 152 -856
rect 106 -1244 112 -868
rect 146 -1244 152 -868
rect 106 -1256 152 -1244
rect -96 -1303 96 -1297
rect -96 -1337 -84 -1303
rect 84 -1337 96 -1303
rect -96 -1343 96 -1337
rect -152 -1396 -106 -1384
rect -152 -1772 -146 -1396
rect -112 -1772 -106 -1396
rect -152 -1784 -106 -1772
rect 106 -1396 152 -1384
rect 106 -1772 112 -1396
rect 146 -1772 152 -1396
rect 106 -1784 152 -1772
rect -96 -1831 96 -1825
rect -96 -1865 -84 -1831
rect 84 -1865 96 -1831
rect -96 -1871 96 -1865
rect -152 -1924 -106 -1912
rect -152 -2300 -146 -1924
rect -112 -2300 -106 -1924
rect -152 -2312 -106 -2300
rect 106 -1924 152 -1912
rect 106 -2300 112 -1924
rect 146 -2300 152 -1924
rect 106 -2312 152 -2300
rect -96 -2359 96 -2353
rect -96 -2393 -84 -2359
rect 84 -2393 96 -2359
rect -96 -2399 96 -2393
rect -152 -2452 -106 -2440
rect -152 -2828 -146 -2452
rect -112 -2828 -106 -2452
rect -152 -2840 -106 -2828
rect 106 -2452 152 -2440
rect 106 -2828 112 -2452
rect 146 -2828 152 -2452
rect 106 -2840 152 -2828
rect -96 -2887 96 -2881
rect -96 -2921 -84 -2887
rect 84 -2921 96 -2887
rect -96 -2927 96 -2921
rect -152 -2980 -106 -2968
rect -152 -3356 -146 -2980
rect -112 -3356 -106 -2980
rect -152 -3368 -106 -3356
rect 106 -2980 152 -2968
rect 106 -3356 112 -2980
rect 146 -3356 152 -2980
rect 106 -3368 152 -3356
rect -96 -3415 96 -3409
rect -96 -3449 -84 -3415
rect 84 -3449 96 -3415
rect -96 -3455 96 -3449
rect -152 -3508 -106 -3496
rect -152 -3884 -146 -3508
rect -112 -3884 -106 -3508
rect -152 -3896 -106 -3884
rect 106 -3508 152 -3496
rect 106 -3884 112 -3508
rect 146 -3884 152 -3508
rect 106 -3896 152 -3884
rect -96 -3943 96 -3937
rect -96 -3977 -84 -3943
rect 84 -3977 96 -3943
rect -96 -3983 96 -3977
<< properties >>
string FIXED_BBOX -263 -4098 263 4098
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 1 m 15 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
